module textFlashTop(

);

// Data is stored in Flash as a binary map of a character
// Example: The following would be a low resolution map of the letter I
//
// 1111111111
// 0000110000
// 0000110000
// 0000110000
// 0000110000
// 1111111111
//
//
// The goal is to have high resolution maps for multiple fonts


// Use caching to improve average memory access time

endmodule
// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 18.0.0 Build 614 04/24/2018 SJ Lite Edition"

// DATE "02/04/2020 21:26:41"

// 
// Device: Altera EP4CE22F17C6 Package FBGA256
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module flashLoader (
	\dut_asmiblock~ALTERA_DCLK ,
	\dut_asmiblock~ALTERA_SCE ,
	\dut_asmiblock~ALTERA_SDO ,
	\dut_asmiblock~ALTERA_DATA0 ,
	avl_csr_address,
	avl_csr_read,
	avl_csr_readdata,
	avl_csr_write,
	avl_csr_writedata,
	avl_csr_waitrequest,
	avl_csr_readdatavalid,
	avl_mem_write,
	avl_mem_burstcount,
	avl_mem_waitrequest,
	avl_mem_read,
	avl_mem_address,
	avl_mem_writedata,
	avl_mem_readdata,
	avl_mem_readdatavalid,
	avl_mem_byteenable,
	clk_clk,
	reset_reset)/* synthesis synthesis_greybox=0 */;
output 	\dut_asmiblock~ALTERA_DCLK ;
output 	\dut_asmiblock~ALTERA_SCE ;
output 	\dut_asmiblock~ALTERA_SDO ;
input 	\dut_asmiblock~ALTERA_DATA0 ;
input 	[5:0] avl_csr_address;
input 	avl_csr_read;
output 	[31:0] avl_csr_readdata;
input 	avl_csr_write;
input 	[31:0] avl_csr_writedata;
output 	avl_csr_waitrequest;
output 	avl_csr_readdatavalid;
input 	avl_mem_write;
input 	[6:0] avl_mem_burstcount;
output 	avl_mem_waitrequest;
input 	avl_mem_read;
input 	[20:0] avl_mem_address;
input 	[31:0] avl_mem_writedata;
output 	[31:0] avl_mem_readdata;
output 	avl_mem_readdatavalid;
input 	[3:0] avl_mem_byteenable;
input 	clk_clk;
input 	reset_reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[0]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[1]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[2]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[3]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[4]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[5]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[6]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[7]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[8]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[9]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[10]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[11]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[12]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[13]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[14]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[15]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[16]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[17]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[18]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[19]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[20]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[21]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[22]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[23]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[24]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[25]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[26]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[27]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[28]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[29]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[30]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[31]~q ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|csr_waitrequest~combout ;
wire \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddatavalid_local~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_waitrequest~0_combout ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[0]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[1]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[2]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[3]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[4]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[5]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[6]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[7]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[8]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[9]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[10]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[11]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[12]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[13]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[14]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[15]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[16]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[17]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[18]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[19]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[20]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[21]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[22]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[23]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[24]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[25]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[26]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[27]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[28]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[29]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[30]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[31]~q ;
wire \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddatavalid~q ;
wire \intel_generic_serial_flash_interface_top_0|qspi_inf_inst|flash_clk_reg~q ;
wire \intel_generic_serial_flash_interface_top_0|qspi_inf_inst|oe_reg~q ;
wire \intel_generic_serial_flash_interface_top_0|qspi_inf_inst|ncs_reg[0]~q ;
wire \intel_generic_serial_flash_interface_top_0|qspi_inf_inst|flash_data_out_reg[0]~q ;
wire \avl_csr_address[1]~input_o ;
wire \avl_csr_address[0]~input_o ;
wire \avl_csr_address[2]~input_o ;
wire \avl_csr_address[3]~input_o ;
wire \avl_csr_read~input_o ;
wire \avl_csr_address[4]~input_o ;
wire \avl_csr_address[5]~input_o ;
wire \clk_clk~input_o ;
wire \avl_csr_write~input_o ;
wire \avl_csr_writedata[0]~input_o ;
wire \avl_csr_writedata[1]~input_o ;
wire \avl_csr_writedata[2]~input_o ;
wire \avl_csr_writedata[3]~input_o ;
wire \avl_csr_writedata[4]~input_o ;
wire \avl_csr_writedata[5]~input_o ;
wire \avl_csr_writedata[6]~input_o ;
wire \avl_csr_writedata[7]~input_o ;
wire \avl_csr_writedata[8]~input_o ;
wire \avl_csr_writedata[9]~input_o ;
wire \avl_csr_writedata[10]~input_o ;
wire \avl_csr_writedata[11]~input_o ;
wire \avl_csr_writedata[12]~input_o ;
wire \avl_csr_writedata[13]~input_o ;
wire \avl_csr_writedata[14]~input_o ;
wire \avl_csr_writedata[15]~input_o ;
wire \avl_csr_writedata[16]~input_o ;
wire \avl_csr_writedata[17]~input_o ;
wire \avl_csr_writedata[18]~input_o ;
wire \avl_csr_writedata[19]~input_o ;
wire \avl_csr_writedata[20]~input_o ;
wire \avl_csr_writedata[21]~input_o ;
wire \avl_csr_writedata[22]~input_o ;
wire \avl_csr_writedata[23]~input_o ;
wire \avl_csr_writedata[24]~input_o ;
wire \avl_csr_writedata[25]~input_o ;
wire \avl_csr_writedata[26]~input_o ;
wire \avl_csr_writedata[27]~input_o ;
wire \avl_csr_writedata[28]~input_o ;
wire \avl_csr_writedata[29]~input_o ;
wire \avl_csr_writedata[30]~input_o ;
wire \avl_csr_writedata[31]~input_o ;
wire \avl_mem_read~input_o ;
wire \avl_mem_burstcount[0]~input_o ;
wire \avl_mem_burstcount[6]~input_o ;
wire \avl_mem_burstcount[2]~input_o ;
wire \avl_mem_burstcount[1]~input_o ;
wire \avl_mem_burstcount[5]~input_o ;
wire \avl_mem_burstcount[4]~input_o ;
wire \avl_mem_burstcount[3]~input_o ;
wire \avl_mem_write~input_o ;
wire \avl_mem_byteenable[0]~input_o ;
wire \avl_mem_byteenable[1]~input_o ;
wire \avl_mem_byteenable[2]~input_o ;
wire \avl_mem_byteenable[3]~input_o ;
wire \reset_reset~input_o ;
wire \avl_mem_writedata[30]~input_o ;
wire \avl_mem_writedata[29]~input_o ;
wire \avl_mem_writedata[28]~input_o ;
wire \avl_mem_writedata[27]~input_o ;
wire \avl_mem_writedata[11]~input_o ;
wire \avl_mem_writedata[18]~input_o ;
wire \avl_mem_writedata[19]~input_o ;
wire \avl_mem_writedata[21]~input_o ;
wire \avl_mem_writedata[20]~input_o ;
wire \avl_mem_writedata[22]~input_o ;
wire \avl_mem_writedata[23]~input_o ;
wire \avl_mem_writedata[24]~input_o ;
wire \avl_mem_writedata[25]~input_o ;
wire \avl_mem_writedata[26]~input_o ;
wire \avl_mem_writedata[10]~input_o ;
wire \avl_mem_writedata[8]~input_o ;
wire \intel_generic_serial_flash_interface_top_0|qspi_inf_inst|dedicated_interface|dut_asmiblock~ALTERA_DATA0input_o ;
wire \avl_mem_writedata[13]~input_o ;
wire \avl_mem_writedata[17]~input_o ;
wire \avl_mem_writedata[16]~input_o ;
wire \avl_mem_writedata[15]~input_o ;
wire \avl_mem_writedata[31]~input_o ;
wire \avl_mem_writedata[14]~input_o ;
wire \avl_mem_writedata[9]~input_o ;
wire \avl_mem_address[6]~input_o ;
wire \avl_mem_address[14]~input_o ;
wire \avl_mem_writedata[0]~input_o ;
wire \avl_mem_address[10]~input_o ;
wire \avl_mem_address[18]~input_o ;
wire \avl_mem_address[2]~input_o ;
wire \avl_mem_writedata[4]~input_o ;
wire \avl_mem_writedata[12]~input_o ;
wire \avl_mem_address[8]~input_o ;
wire \avl_mem_address[16]~input_o ;
wire \avl_mem_address[0]~input_o ;
wire \avl_mem_writedata[2]~input_o ;
wire \avl_mem_address[15]~input_o ;
wire \avl_mem_address[7]~input_o ;
wire \avl_mem_writedata[1]~input_o ;
wire \avl_mem_address[17]~input_o ;
wire \avl_mem_address[9]~input_o ;
wire \avl_mem_address[1]~input_o ;
wire \avl_mem_writedata[3]~input_o ;
wire \avl_mem_address[19]~input_o ;
wire \avl_mem_address[11]~input_o ;
wire \avl_mem_address[3]~input_o ;
wire \avl_mem_writedata[5]~input_o ;
wire \avl_mem_address[12]~input_o ;
wire \avl_mem_address[20]~input_o ;
wire \avl_mem_address[4]~input_o ;
wire \avl_mem_writedata[6]~input_o ;
wire \avl_mem_address[13]~input_o ;
wire \avl_mem_address[5]~input_o ;
wire \avl_mem_writedata[7]~input_o ;


flashLoader_flashLoader_intel_generic_serial_flash_interface_top_0 intel_generic_serial_flash_interface_top_0(
	.avl_rddata_local_0(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[0]~q ),
	.avl_rddata_local_1(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[1]~q ),
	.avl_rddata_local_2(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[2]~q ),
	.avl_rddata_local_3(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[3]~q ),
	.avl_rddata_local_4(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[4]~q ),
	.avl_rddata_local_5(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[5]~q ),
	.avl_rddata_local_6(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[6]~q ),
	.avl_rddata_local_7(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[7]~q ),
	.avl_rddata_local_8(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[8]~q ),
	.avl_rddata_local_9(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[9]~q ),
	.avl_rddata_local_10(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[10]~q ),
	.avl_rddata_local_11(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[11]~q ),
	.avl_rddata_local_12(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[12]~q ),
	.avl_rddata_local_13(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[13]~q ),
	.avl_rddata_local_14(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[14]~q ),
	.avl_rddata_local_15(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[15]~q ),
	.avl_rddata_local_16(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[16]~q ),
	.avl_rddata_local_17(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[17]~q ),
	.avl_rddata_local_18(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[18]~q ),
	.avl_rddata_local_19(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[19]~q ),
	.avl_rddata_local_20(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[20]~q ),
	.avl_rddata_local_21(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[21]~q ),
	.avl_rddata_local_22(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[22]~q ),
	.avl_rddata_local_23(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[23]~q ),
	.avl_rddata_local_24(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[24]~q ),
	.avl_rddata_local_25(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[25]~q ),
	.avl_rddata_local_26(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[26]~q ),
	.avl_rddata_local_27(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[27]~q ),
	.avl_rddata_local_28(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[28]~q ),
	.avl_rddata_local_29(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[29]~q ),
	.avl_rddata_local_30(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[30]~q ),
	.avl_rddata_local_31(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[31]~q ),
	.csr_waitrequest(\intel_generic_serial_flash_interface_top_0|csr_controller|csr_waitrequest~combout ),
	.avl_rddatavalid_local(\intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddatavalid_local~q ),
	.mem_waitrequest(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_waitrequest~0_combout ),
	.mem_rddata_0(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[0]~q ),
	.mem_rddata_1(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[1]~q ),
	.mem_rddata_2(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[2]~q ),
	.mem_rddata_3(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[3]~q ),
	.mem_rddata_4(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[4]~q ),
	.mem_rddata_5(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[5]~q ),
	.mem_rddata_6(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[6]~q ),
	.mem_rddata_7(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[7]~q ),
	.mem_rddata_8(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[8]~q ),
	.mem_rddata_9(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[9]~q ),
	.mem_rddata_10(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[10]~q ),
	.mem_rddata_11(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[11]~q ),
	.mem_rddata_12(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[12]~q ),
	.mem_rddata_13(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[13]~q ),
	.mem_rddata_14(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[14]~q ),
	.mem_rddata_15(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[15]~q ),
	.mem_rddata_16(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[16]~q ),
	.mem_rddata_17(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[17]~q ),
	.mem_rddata_18(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[18]~q ),
	.mem_rddata_19(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[19]~q ),
	.mem_rddata_20(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[20]~q ),
	.mem_rddata_21(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[21]~q ),
	.mem_rddata_22(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[22]~q ),
	.mem_rddata_23(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[23]~q ),
	.mem_rddata_24(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[24]~q ),
	.mem_rddata_25(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[25]~q ),
	.mem_rddata_26(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[26]~q ),
	.mem_rddata_27(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[27]~q ),
	.mem_rddata_28(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[28]~q ),
	.mem_rddata_29(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[29]~q ),
	.mem_rddata_30(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[30]~q ),
	.mem_rddata_31(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[31]~q ),
	.mem_rddatavalid(\intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddatavalid~q ),
	.flash_clk_reg(\intel_generic_serial_flash_interface_top_0|qspi_inf_inst|flash_clk_reg~q ),
	.oe_reg(\intel_generic_serial_flash_interface_top_0|qspi_inf_inst|oe_reg~q ),
	.ncs_reg_0(\intel_generic_serial_flash_interface_top_0|qspi_inf_inst|ncs_reg[0]~q ),
	.flash_data_out_reg_0(\intel_generic_serial_flash_interface_top_0|qspi_inf_inst|flash_data_out_reg[0]~q ),
	.avl_csr_address_1(\avl_csr_address[1]~input_o ),
	.avl_csr_address_0(\avl_csr_address[0]~input_o ),
	.avl_csr_address_2(\avl_csr_address[2]~input_o ),
	.avl_csr_address_3(\avl_csr_address[3]~input_o ),
	.avl_csr_read(\avl_csr_read~input_o ),
	.avl_csr_address_4(\avl_csr_address[4]~input_o ),
	.avl_csr_address_5(\avl_csr_address[5]~input_o ),
	.clk_clk(\clk_clk~input_o ),
	.avl_csr_write(\avl_csr_write~input_o ),
	.avl_csr_writedata_0(\avl_csr_writedata[0]~input_o ),
	.avl_csr_writedata_1(\avl_csr_writedata[1]~input_o ),
	.avl_csr_writedata_2(\avl_csr_writedata[2]~input_o ),
	.avl_csr_writedata_3(\avl_csr_writedata[3]~input_o ),
	.avl_csr_writedata_4(\avl_csr_writedata[4]~input_o ),
	.avl_csr_writedata_5(\avl_csr_writedata[5]~input_o ),
	.avl_csr_writedata_6(\avl_csr_writedata[6]~input_o ),
	.avl_csr_writedata_7(\avl_csr_writedata[7]~input_o ),
	.avl_csr_writedata_8(\avl_csr_writedata[8]~input_o ),
	.avl_csr_writedata_9(\avl_csr_writedata[9]~input_o ),
	.avl_csr_writedata_10(\avl_csr_writedata[10]~input_o ),
	.avl_csr_writedata_11(\avl_csr_writedata[11]~input_o ),
	.avl_csr_writedata_12(\avl_csr_writedata[12]~input_o ),
	.avl_csr_writedata_13(\avl_csr_writedata[13]~input_o ),
	.avl_csr_writedata_14(\avl_csr_writedata[14]~input_o ),
	.avl_csr_writedata_15(\avl_csr_writedata[15]~input_o ),
	.avl_csr_writedata_16(\avl_csr_writedata[16]~input_o ),
	.avl_csr_writedata_17(\avl_csr_writedata[17]~input_o ),
	.avl_csr_writedata_18(\avl_csr_writedata[18]~input_o ),
	.avl_csr_writedata_19(\avl_csr_writedata[19]~input_o ),
	.avl_csr_writedata_20(\avl_csr_writedata[20]~input_o ),
	.avl_csr_writedata_21(\avl_csr_writedata[21]~input_o ),
	.avl_csr_writedata_22(\avl_csr_writedata[22]~input_o ),
	.avl_csr_writedata_23(\avl_csr_writedata[23]~input_o ),
	.avl_csr_writedata_24(\avl_csr_writedata[24]~input_o ),
	.avl_csr_writedata_25(\avl_csr_writedata[25]~input_o ),
	.avl_csr_writedata_26(\avl_csr_writedata[26]~input_o ),
	.avl_csr_writedata_27(\avl_csr_writedata[27]~input_o ),
	.avl_csr_writedata_28(\avl_csr_writedata[28]~input_o ),
	.avl_csr_writedata_29(\avl_csr_writedata[29]~input_o ),
	.avl_csr_writedata_30(\avl_csr_writedata[30]~input_o ),
	.avl_csr_writedata_31(\avl_csr_writedata[31]~input_o ),
	.avl_mem_read(\avl_mem_read~input_o ),
	.avl_mem_burstcount_0(\avl_mem_burstcount[0]~input_o ),
	.avl_mem_burstcount_6(\avl_mem_burstcount[6]~input_o ),
	.avl_mem_burstcount_2(\avl_mem_burstcount[2]~input_o ),
	.avl_mem_burstcount_1(\avl_mem_burstcount[1]~input_o ),
	.avl_mem_burstcount_5(\avl_mem_burstcount[5]~input_o ),
	.avl_mem_burstcount_4(\avl_mem_burstcount[4]~input_o ),
	.avl_mem_burstcount_3(\avl_mem_burstcount[3]~input_o ),
	.avl_mem_write(\avl_mem_write~input_o ),
	.avl_mem_byteenable_0(\avl_mem_byteenable[0]~input_o ),
	.avl_mem_byteenable_1(\avl_mem_byteenable[1]~input_o ),
	.avl_mem_byteenable_2(\avl_mem_byteenable[2]~input_o ),
	.avl_mem_byteenable_3(\avl_mem_byteenable[3]~input_o ),
	.reset_reset(\reset_reset~input_o ),
	.avl_mem_writedata_30(\avl_mem_writedata[30]~input_o ),
	.avl_mem_writedata_29(\avl_mem_writedata[29]~input_o ),
	.avl_mem_writedata_28(\avl_mem_writedata[28]~input_o ),
	.avl_mem_writedata_27(\avl_mem_writedata[27]~input_o ),
	.avl_mem_writedata_11(\avl_mem_writedata[11]~input_o ),
	.avl_mem_writedata_18(\avl_mem_writedata[18]~input_o ),
	.avl_mem_writedata_19(\avl_mem_writedata[19]~input_o ),
	.avl_mem_writedata_21(\avl_mem_writedata[21]~input_o ),
	.avl_mem_writedata_20(\avl_mem_writedata[20]~input_o ),
	.avl_mem_writedata_22(\avl_mem_writedata[22]~input_o ),
	.avl_mem_writedata_23(\avl_mem_writedata[23]~input_o ),
	.avl_mem_writedata_24(\avl_mem_writedata[24]~input_o ),
	.avl_mem_writedata_25(\avl_mem_writedata[25]~input_o ),
	.avl_mem_writedata_26(\avl_mem_writedata[26]~input_o ),
	.avl_mem_writedata_10(\avl_mem_writedata[10]~input_o ),
	.avl_mem_writedata_8(\avl_mem_writedata[8]~input_o ),
	.dut_asmiblock(\intel_generic_serial_flash_interface_top_0|qspi_inf_inst|dedicated_interface|dut_asmiblock~ALTERA_DATA0input_o ),
	.avl_mem_writedata_13(\avl_mem_writedata[13]~input_o ),
	.avl_mem_writedata_17(\avl_mem_writedata[17]~input_o ),
	.avl_mem_writedata_16(\avl_mem_writedata[16]~input_o ),
	.avl_mem_writedata_15(\avl_mem_writedata[15]~input_o ),
	.avl_mem_writedata_31(\avl_mem_writedata[31]~input_o ),
	.avl_mem_writedata_14(\avl_mem_writedata[14]~input_o ),
	.avl_mem_writedata_9(\avl_mem_writedata[9]~input_o ),
	.avl_mem_address_6(\avl_mem_address[6]~input_o ),
	.avl_mem_address_14(\avl_mem_address[14]~input_o ),
	.avl_mem_writedata_0(\avl_mem_writedata[0]~input_o ),
	.avl_mem_address_10(\avl_mem_address[10]~input_o ),
	.avl_mem_address_18(\avl_mem_address[18]~input_o ),
	.avl_mem_address_2(\avl_mem_address[2]~input_o ),
	.avl_mem_writedata_4(\avl_mem_writedata[4]~input_o ),
	.avl_mem_writedata_12(\avl_mem_writedata[12]~input_o ),
	.avl_mem_address_8(\avl_mem_address[8]~input_o ),
	.avl_mem_address_16(\avl_mem_address[16]~input_o ),
	.avl_mem_address_0(\avl_mem_address[0]~input_o ),
	.avl_mem_writedata_2(\avl_mem_writedata[2]~input_o ),
	.avl_mem_address_15(\avl_mem_address[15]~input_o ),
	.avl_mem_address_7(\avl_mem_address[7]~input_o ),
	.avl_mem_writedata_1(\avl_mem_writedata[1]~input_o ),
	.avl_mem_address_17(\avl_mem_address[17]~input_o ),
	.avl_mem_address_9(\avl_mem_address[9]~input_o ),
	.avl_mem_address_1(\avl_mem_address[1]~input_o ),
	.avl_mem_writedata_3(\avl_mem_writedata[3]~input_o ),
	.avl_mem_address_19(\avl_mem_address[19]~input_o ),
	.avl_mem_address_11(\avl_mem_address[11]~input_o ),
	.avl_mem_address_3(\avl_mem_address[3]~input_o ),
	.avl_mem_writedata_5(\avl_mem_writedata[5]~input_o ),
	.avl_mem_address_12(\avl_mem_address[12]~input_o ),
	.avl_mem_address_20(\avl_mem_address[20]~input_o ),
	.avl_mem_address_4(\avl_mem_address[4]~input_o ),
	.avl_mem_writedata_6(\avl_mem_writedata[6]~input_o ),
	.avl_mem_address_13(\avl_mem_address[13]~input_o ),
	.avl_mem_address_5(\avl_mem_address[5]~input_o ),
	.avl_mem_writedata_7(\avl_mem_writedata[7]~input_o ));

assign \avl_csr_address[1]~input_o  = avl_csr_address[1];

assign \avl_csr_address[0]~input_o  = avl_csr_address[0];

assign \avl_csr_address[2]~input_o  = avl_csr_address[2];

assign \avl_csr_address[3]~input_o  = avl_csr_address[3];

assign \avl_csr_read~input_o  = avl_csr_read;

assign \avl_csr_address[4]~input_o  = avl_csr_address[4];

assign \avl_csr_address[5]~input_o  = avl_csr_address[5];

assign \clk_clk~input_o  = clk_clk;

assign \avl_csr_write~input_o  = avl_csr_write;

assign \avl_csr_writedata[0]~input_o  = avl_csr_writedata[0];

assign \avl_csr_writedata[1]~input_o  = avl_csr_writedata[1];

assign \avl_csr_writedata[2]~input_o  = avl_csr_writedata[2];

assign \avl_csr_writedata[3]~input_o  = avl_csr_writedata[3];

assign \avl_csr_writedata[4]~input_o  = avl_csr_writedata[4];

assign \avl_csr_writedata[5]~input_o  = avl_csr_writedata[5];

assign \avl_csr_writedata[6]~input_o  = avl_csr_writedata[6];

assign \avl_csr_writedata[7]~input_o  = avl_csr_writedata[7];

assign \avl_csr_writedata[8]~input_o  = avl_csr_writedata[8];

assign \avl_csr_writedata[9]~input_o  = avl_csr_writedata[9];

assign \avl_csr_writedata[10]~input_o  = avl_csr_writedata[10];

assign \avl_csr_writedata[11]~input_o  = avl_csr_writedata[11];

assign \avl_csr_writedata[12]~input_o  = avl_csr_writedata[12];

assign \avl_csr_writedata[13]~input_o  = avl_csr_writedata[13];

assign \avl_csr_writedata[14]~input_o  = avl_csr_writedata[14];

assign \avl_csr_writedata[15]~input_o  = avl_csr_writedata[15];

assign \avl_csr_writedata[16]~input_o  = avl_csr_writedata[16];

assign \avl_csr_writedata[17]~input_o  = avl_csr_writedata[17];

assign \avl_csr_writedata[18]~input_o  = avl_csr_writedata[18];

assign \avl_csr_writedata[19]~input_o  = avl_csr_writedata[19];

assign \avl_csr_writedata[20]~input_o  = avl_csr_writedata[20];

assign \avl_csr_writedata[21]~input_o  = avl_csr_writedata[21];

assign \avl_csr_writedata[22]~input_o  = avl_csr_writedata[22];

assign \avl_csr_writedata[23]~input_o  = avl_csr_writedata[23];

assign \avl_csr_writedata[24]~input_o  = avl_csr_writedata[24];

assign \avl_csr_writedata[25]~input_o  = avl_csr_writedata[25];

assign \avl_csr_writedata[26]~input_o  = avl_csr_writedata[26];

assign \avl_csr_writedata[27]~input_o  = avl_csr_writedata[27];

assign \avl_csr_writedata[28]~input_o  = avl_csr_writedata[28];

assign \avl_csr_writedata[29]~input_o  = avl_csr_writedata[29];

assign \avl_csr_writedata[30]~input_o  = avl_csr_writedata[30];

assign \avl_csr_writedata[31]~input_o  = avl_csr_writedata[31];

assign \avl_mem_read~input_o  = avl_mem_read;

assign \avl_mem_burstcount[0]~input_o  = avl_mem_burstcount[0];

assign \avl_mem_burstcount[6]~input_o  = avl_mem_burstcount[6];

assign \avl_mem_burstcount[2]~input_o  = avl_mem_burstcount[2];

assign \avl_mem_burstcount[1]~input_o  = avl_mem_burstcount[1];

assign \avl_mem_burstcount[5]~input_o  = avl_mem_burstcount[5];

assign \avl_mem_burstcount[4]~input_o  = avl_mem_burstcount[4];

assign \avl_mem_burstcount[3]~input_o  = avl_mem_burstcount[3];

assign \avl_mem_write~input_o  = avl_mem_write;

assign \avl_mem_byteenable[0]~input_o  = avl_mem_byteenable[0];

assign \avl_mem_byteenable[1]~input_o  = avl_mem_byteenable[1];

assign \avl_mem_byteenable[2]~input_o  = avl_mem_byteenable[2];

assign \avl_mem_byteenable[3]~input_o  = avl_mem_byteenable[3];

assign \reset_reset~input_o  = reset_reset;

assign \avl_mem_writedata[30]~input_o  = avl_mem_writedata[30];

assign \avl_mem_writedata[29]~input_o  = avl_mem_writedata[29];

assign \avl_mem_writedata[28]~input_o  = avl_mem_writedata[28];

assign \avl_mem_writedata[27]~input_o  = avl_mem_writedata[27];

assign \avl_mem_writedata[11]~input_o  = avl_mem_writedata[11];

assign \avl_mem_writedata[18]~input_o  = avl_mem_writedata[18];

assign \avl_mem_writedata[19]~input_o  = avl_mem_writedata[19];

assign \avl_mem_writedata[21]~input_o  = avl_mem_writedata[21];

assign \avl_mem_writedata[20]~input_o  = avl_mem_writedata[20];

assign \avl_mem_writedata[22]~input_o  = avl_mem_writedata[22];

assign \avl_mem_writedata[23]~input_o  = avl_mem_writedata[23];

assign \avl_mem_writedata[24]~input_o  = avl_mem_writedata[24];

assign \avl_mem_writedata[25]~input_o  = avl_mem_writedata[25];

assign \avl_mem_writedata[26]~input_o  = avl_mem_writedata[26];

assign \avl_mem_writedata[10]~input_o  = avl_mem_writedata[10];

assign \avl_mem_writedata[8]~input_o  = avl_mem_writedata[8];

assign \intel_generic_serial_flash_interface_top_0|qspi_inf_inst|dedicated_interface|dut_asmiblock~ALTERA_DATA0input_o  = \dut_asmiblock~ALTERA_DATA0 ;

assign \avl_mem_writedata[13]~input_o  = avl_mem_writedata[13];

assign \avl_mem_writedata[17]~input_o  = avl_mem_writedata[17];

assign \avl_mem_writedata[16]~input_o  = avl_mem_writedata[16];

assign \avl_mem_writedata[15]~input_o  = avl_mem_writedata[15];

assign \avl_mem_writedata[31]~input_o  = avl_mem_writedata[31];

assign \avl_mem_writedata[14]~input_o  = avl_mem_writedata[14];

assign \avl_mem_writedata[9]~input_o  = avl_mem_writedata[9];

assign \avl_mem_address[6]~input_o  = avl_mem_address[6];

assign \avl_mem_address[14]~input_o  = avl_mem_address[14];

assign \avl_mem_writedata[0]~input_o  = avl_mem_writedata[0];

assign \avl_mem_address[10]~input_o  = avl_mem_address[10];

assign \avl_mem_address[18]~input_o  = avl_mem_address[18];

assign \avl_mem_address[2]~input_o  = avl_mem_address[2];

assign \avl_mem_writedata[4]~input_o  = avl_mem_writedata[4];

assign \avl_mem_writedata[12]~input_o  = avl_mem_writedata[12];

assign \avl_mem_address[8]~input_o  = avl_mem_address[8];

assign \avl_mem_address[16]~input_o  = avl_mem_address[16];

assign \avl_mem_address[0]~input_o  = avl_mem_address[0];

assign \avl_mem_writedata[2]~input_o  = avl_mem_writedata[2];

assign \avl_mem_address[15]~input_o  = avl_mem_address[15];

assign \avl_mem_address[7]~input_o  = avl_mem_address[7];

assign \avl_mem_writedata[1]~input_o  = avl_mem_writedata[1];

assign \avl_mem_address[17]~input_o  = avl_mem_address[17];

assign \avl_mem_address[9]~input_o  = avl_mem_address[9];

assign \avl_mem_address[1]~input_o  = avl_mem_address[1];

assign \avl_mem_writedata[3]~input_o  = avl_mem_writedata[3];

assign \avl_mem_address[19]~input_o  = avl_mem_address[19];

assign \avl_mem_address[11]~input_o  = avl_mem_address[11];

assign \avl_mem_address[3]~input_o  = avl_mem_address[3];

assign \avl_mem_writedata[5]~input_o  = avl_mem_writedata[5];

assign \avl_mem_address[12]~input_o  = avl_mem_address[12];

assign \avl_mem_address[20]~input_o  = avl_mem_address[20];

assign \avl_mem_address[4]~input_o  = avl_mem_address[4];

assign \avl_mem_writedata[6]~input_o  = avl_mem_writedata[6];

assign \avl_mem_address[13]~input_o  = avl_mem_address[13];

assign \avl_mem_address[5]~input_o  = avl_mem_address[5];

assign \avl_mem_writedata[7]~input_o  = avl_mem_writedata[7];

cycloneive_io_obuf \intel_generic_serial_flash_interface_top_0|qspi_inf_inst|dedicated_interface|dut_asmiblock~ALTERA_DCLK_OBUF (
	.i(\intel_generic_serial_flash_interface_top_0|qspi_inf_inst|flash_clk_reg~q ),
	.oe(!\intel_generic_serial_flash_interface_top_0|qspi_inf_inst|oe_reg~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(\dut_asmiblock~ALTERA_DCLK ),
	.obar());
defparam \intel_generic_serial_flash_interface_top_0|qspi_inf_inst|dedicated_interface|dut_asmiblock~ALTERA_DCLK_OBUF .bus_hold = "false";
defparam \intel_generic_serial_flash_interface_top_0|qspi_inf_inst|dedicated_interface|dut_asmiblock~ALTERA_DCLK_OBUF .open_drain_output = "false";

cycloneive_io_obuf \intel_generic_serial_flash_interface_top_0|qspi_inf_inst|dedicated_interface|dut_asmiblock~ALTERA_SCE_OBUF (
	.i(!\intel_generic_serial_flash_interface_top_0|qspi_inf_inst|ncs_reg[0]~q ),
	.oe(!\intel_generic_serial_flash_interface_top_0|qspi_inf_inst|oe_reg~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(\dut_asmiblock~ALTERA_SCE ),
	.obar());
defparam \intel_generic_serial_flash_interface_top_0|qspi_inf_inst|dedicated_interface|dut_asmiblock~ALTERA_SCE_OBUF .bus_hold = "false";
defparam \intel_generic_serial_flash_interface_top_0|qspi_inf_inst|dedicated_interface|dut_asmiblock~ALTERA_SCE_OBUF .open_drain_output = "false";

cycloneive_io_obuf \intel_generic_serial_flash_interface_top_0|qspi_inf_inst|dedicated_interface|dut_asmiblock~ALTERA_SDO_OBUF (
	.i(\intel_generic_serial_flash_interface_top_0|qspi_inf_inst|flash_data_out_reg[0]~q ),
	.oe(!\intel_generic_serial_flash_interface_top_0|qspi_inf_inst|oe_reg~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(\dut_asmiblock~ALTERA_SDO ),
	.obar());
defparam \intel_generic_serial_flash_interface_top_0|qspi_inf_inst|dedicated_interface|dut_asmiblock~ALTERA_SDO_OBUF .bus_hold = "false";
defparam \intel_generic_serial_flash_interface_top_0|qspi_inf_inst|dedicated_interface|dut_asmiblock~ALTERA_SDO_OBUF .open_drain_output = "false";

assign avl_csr_readdata[0] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[0]~q ;

assign avl_csr_readdata[1] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[1]~q ;

assign avl_csr_readdata[2] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[2]~q ;

assign avl_csr_readdata[3] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[3]~q ;

assign avl_csr_readdata[4] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[4]~q ;

assign avl_csr_readdata[5] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[5]~q ;

assign avl_csr_readdata[6] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[6]~q ;

assign avl_csr_readdata[7] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[7]~q ;

assign avl_csr_readdata[8] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[8]~q ;

assign avl_csr_readdata[9] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[9]~q ;

assign avl_csr_readdata[10] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[10]~q ;

assign avl_csr_readdata[11] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[11]~q ;

assign avl_csr_readdata[12] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[12]~q ;

assign avl_csr_readdata[13] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[13]~q ;

assign avl_csr_readdata[14] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[14]~q ;

assign avl_csr_readdata[15] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[15]~q ;

assign avl_csr_readdata[16] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[16]~q ;

assign avl_csr_readdata[17] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[17]~q ;

assign avl_csr_readdata[18] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[18]~q ;

assign avl_csr_readdata[19] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[19]~q ;

assign avl_csr_readdata[20] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[20]~q ;

assign avl_csr_readdata[21] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[21]~q ;

assign avl_csr_readdata[22] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[22]~q ;

assign avl_csr_readdata[23] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[23]~q ;

assign avl_csr_readdata[24] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[24]~q ;

assign avl_csr_readdata[25] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[25]~q ;

assign avl_csr_readdata[26] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[26]~q ;

assign avl_csr_readdata[27] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[27]~q ;

assign avl_csr_readdata[28] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[28]~q ;

assign avl_csr_readdata[29] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[29]~q ;

assign avl_csr_readdata[30] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[30]~q ;

assign avl_csr_readdata[31] = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddata_local[31]~q ;

assign avl_csr_waitrequest = \intel_generic_serial_flash_interface_top_0|csr_controller|csr_waitrequest~combout ;

assign avl_csr_readdatavalid = \intel_generic_serial_flash_interface_top_0|csr_controller|avl_rddatavalid_local~q ;

assign avl_mem_waitrequest = ~ \intel_generic_serial_flash_interface_top_0|xip_controller|mem_waitrequest~0_combout ;

assign avl_mem_readdata[0] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[0]~q ;

assign avl_mem_readdata[1] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[1]~q ;

assign avl_mem_readdata[2] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[2]~q ;

assign avl_mem_readdata[3] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[3]~q ;

assign avl_mem_readdata[4] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[4]~q ;

assign avl_mem_readdata[5] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[5]~q ;

assign avl_mem_readdata[6] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[6]~q ;

assign avl_mem_readdata[7] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[7]~q ;

assign avl_mem_readdata[8] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[8]~q ;

assign avl_mem_readdata[9] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[9]~q ;

assign avl_mem_readdata[10] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[10]~q ;

assign avl_mem_readdata[11] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[11]~q ;

assign avl_mem_readdata[12] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[12]~q ;

assign avl_mem_readdata[13] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[13]~q ;

assign avl_mem_readdata[14] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[14]~q ;

assign avl_mem_readdata[15] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[15]~q ;

assign avl_mem_readdata[16] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[16]~q ;

assign avl_mem_readdata[17] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[17]~q ;

assign avl_mem_readdata[18] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[18]~q ;

assign avl_mem_readdata[19] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[19]~q ;

assign avl_mem_readdata[20] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[20]~q ;

assign avl_mem_readdata[21] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[21]~q ;

assign avl_mem_readdata[22] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[22]~q ;

assign avl_mem_readdata[23] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[23]~q ;

assign avl_mem_readdata[24] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[24]~q ;

assign avl_mem_readdata[25] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[25]~q ;

assign avl_mem_readdata[26] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[26]~q ;

assign avl_mem_readdata[27] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[27]~q ;

assign avl_mem_readdata[28] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[28]~q ;

assign avl_mem_readdata[29] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[29]~q ;

assign avl_mem_readdata[30] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[30]~q ;

assign avl_mem_readdata[31] = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddata[31]~q ;

assign avl_mem_readdatavalid = \intel_generic_serial_flash_interface_top_0|xip_controller|mem_rddatavalid~q ;

endmodule

module flashLoader_flashLoader_intel_generic_serial_flash_interface_top_0 (
	avl_rddata_local_0,
	avl_rddata_local_1,
	avl_rddata_local_2,
	avl_rddata_local_3,
	avl_rddata_local_4,
	avl_rddata_local_5,
	avl_rddata_local_6,
	avl_rddata_local_7,
	avl_rddata_local_8,
	avl_rddata_local_9,
	avl_rddata_local_10,
	avl_rddata_local_11,
	avl_rddata_local_12,
	avl_rddata_local_13,
	avl_rddata_local_14,
	avl_rddata_local_15,
	avl_rddata_local_16,
	avl_rddata_local_17,
	avl_rddata_local_18,
	avl_rddata_local_19,
	avl_rddata_local_20,
	avl_rddata_local_21,
	avl_rddata_local_22,
	avl_rddata_local_23,
	avl_rddata_local_24,
	avl_rddata_local_25,
	avl_rddata_local_26,
	avl_rddata_local_27,
	avl_rddata_local_28,
	avl_rddata_local_29,
	avl_rddata_local_30,
	avl_rddata_local_31,
	csr_waitrequest,
	avl_rddatavalid_local,
	mem_waitrequest,
	mem_rddata_0,
	mem_rddata_1,
	mem_rddata_2,
	mem_rddata_3,
	mem_rddata_4,
	mem_rddata_5,
	mem_rddata_6,
	mem_rddata_7,
	mem_rddata_8,
	mem_rddata_9,
	mem_rddata_10,
	mem_rddata_11,
	mem_rddata_12,
	mem_rddata_13,
	mem_rddata_14,
	mem_rddata_15,
	mem_rddata_16,
	mem_rddata_17,
	mem_rddata_18,
	mem_rddata_19,
	mem_rddata_20,
	mem_rddata_21,
	mem_rddata_22,
	mem_rddata_23,
	mem_rddata_24,
	mem_rddata_25,
	mem_rddata_26,
	mem_rddata_27,
	mem_rddata_28,
	mem_rddata_29,
	mem_rddata_30,
	mem_rddata_31,
	mem_rddatavalid,
	flash_clk_reg,
	oe_reg,
	ncs_reg_0,
	flash_data_out_reg_0,
	avl_csr_address_1,
	avl_csr_address_0,
	avl_csr_address_2,
	avl_csr_address_3,
	avl_csr_read,
	avl_csr_address_4,
	avl_csr_address_5,
	clk_clk,
	avl_csr_write,
	avl_csr_writedata_0,
	avl_csr_writedata_1,
	avl_csr_writedata_2,
	avl_csr_writedata_3,
	avl_csr_writedata_4,
	avl_csr_writedata_5,
	avl_csr_writedata_6,
	avl_csr_writedata_7,
	avl_csr_writedata_8,
	avl_csr_writedata_9,
	avl_csr_writedata_10,
	avl_csr_writedata_11,
	avl_csr_writedata_12,
	avl_csr_writedata_13,
	avl_csr_writedata_14,
	avl_csr_writedata_15,
	avl_csr_writedata_16,
	avl_csr_writedata_17,
	avl_csr_writedata_18,
	avl_csr_writedata_19,
	avl_csr_writedata_20,
	avl_csr_writedata_21,
	avl_csr_writedata_22,
	avl_csr_writedata_23,
	avl_csr_writedata_24,
	avl_csr_writedata_25,
	avl_csr_writedata_26,
	avl_csr_writedata_27,
	avl_csr_writedata_28,
	avl_csr_writedata_29,
	avl_csr_writedata_30,
	avl_csr_writedata_31,
	avl_mem_read,
	avl_mem_burstcount_0,
	avl_mem_burstcount_6,
	avl_mem_burstcount_2,
	avl_mem_burstcount_1,
	avl_mem_burstcount_5,
	avl_mem_burstcount_4,
	avl_mem_burstcount_3,
	avl_mem_write,
	avl_mem_byteenable_0,
	avl_mem_byteenable_1,
	avl_mem_byteenable_2,
	avl_mem_byteenable_3,
	reset_reset,
	avl_mem_writedata_30,
	avl_mem_writedata_29,
	avl_mem_writedata_28,
	avl_mem_writedata_27,
	avl_mem_writedata_11,
	avl_mem_writedata_18,
	avl_mem_writedata_19,
	avl_mem_writedata_21,
	avl_mem_writedata_20,
	avl_mem_writedata_22,
	avl_mem_writedata_23,
	avl_mem_writedata_24,
	avl_mem_writedata_25,
	avl_mem_writedata_26,
	avl_mem_writedata_10,
	avl_mem_writedata_8,
	dut_asmiblock,
	avl_mem_writedata_13,
	avl_mem_writedata_17,
	avl_mem_writedata_16,
	avl_mem_writedata_15,
	avl_mem_writedata_31,
	avl_mem_writedata_14,
	avl_mem_writedata_9,
	avl_mem_address_6,
	avl_mem_address_14,
	avl_mem_writedata_0,
	avl_mem_address_10,
	avl_mem_address_18,
	avl_mem_address_2,
	avl_mem_writedata_4,
	avl_mem_writedata_12,
	avl_mem_address_8,
	avl_mem_address_16,
	avl_mem_address_0,
	avl_mem_writedata_2,
	avl_mem_address_15,
	avl_mem_address_7,
	avl_mem_writedata_1,
	avl_mem_address_17,
	avl_mem_address_9,
	avl_mem_address_1,
	avl_mem_writedata_3,
	avl_mem_address_19,
	avl_mem_address_11,
	avl_mem_address_3,
	avl_mem_writedata_5,
	avl_mem_address_12,
	avl_mem_address_20,
	avl_mem_address_4,
	avl_mem_writedata_6,
	avl_mem_address_13,
	avl_mem_address_5,
	avl_mem_writedata_7)/* synthesis synthesis_greybox=0 */;
output 	avl_rddata_local_0;
output 	avl_rddata_local_1;
output 	avl_rddata_local_2;
output 	avl_rddata_local_3;
output 	avl_rddata_local_4;
output 	avl_rddata_local_5;
output 	avl_rddata_local_6;
output 	avl_rddata_local_7;
output 	avl_rddata_local_8;
output 	avl_rddata_local_9;
output 	avl_rddata_local_10;
output 	avl_rddata_local_11;
output 	avl_rddata_local_12;
output 	avl_rddata_local_13;
output 	avl_rddata_local_14;
output 	avl_rddata_local_15;
output 	avl_rddata_local_16;
output 	avl_rddata_local_17;
output 	avl_rddata_local_18;
output 	avl_rddata_local_19;
output 	avl_rddata_local_20;
output 	avl_rddata_local_21;
output 	avl_rddata_local_22;
output 	avl_rddata_local_23;
output 	avl_rddata_local_24;
output 	avl_rddata_local_25;
output 	avl_rddata_local_26;
output 	avl_rddata_local_27;
output 	avl_rddata_local_28;
output 	avl_rddata_local_29;
output 	avl_rddata_local_30;
output 	avl_rddata_local_31;
output 	csr_waitrequest;
output 	avl_rddatavalid_local;
output 	mem_waitrequest;
output 	mem_rddata_0;
output 	mem_rddata_1;
output 	mem_rddata_2;
output 	mem_rddata_3;
output 	mem_rddata_4;
output 	mem_rddata_5;
output 	mem_rddata_6;
output 	mem_rddata_7;
output 	mem_rddata_8;
output 	mem_rddata_9;
output 	mem_rddata_10;
output 	mem_rddata_11;
output 	mem_rddata_12;
output 	mem_rddata_13;
output 	mem_rddata_14;
output 	mem_rddata_15;
output 	mem_rddata_16;
output 	mem_rddata_17;
output 	mem_rddata_18;
output 	mem_rddata_19;
output 	mem_rddata_20;
output 	mem_rddata_21;
output 	mem_rddata_22;
output 	mem_rddata_23;
output 	mem_rddata_24;
output 	mem_rddata_25;
output 	mem_rddata_26;
output 	mem_rddata_27;
output 	mem_rddata_28;
output 	mem_rddata_29;
output 	mem_rddata_30;
output 	mem_rddata_31;
output 	mem_rddatavalid;
output 	flash_clk_reg;
output 	oe_reg;
output 	ncs_reg_0;
output 	flash_data_out_reg_0;
input 	avl_csr_address_1;
input 	avl_csr_address_0;
input 	avl_csr_address_2;
input 	avl_csr_address_3;
input 	avl_csr_read;
input 	avl_csr_address_4;
input 	avl_csr_address_5;
input 	clk_clk;
input 	avl_csr_write;
input 	avl_csr_writedata_0;
input 	avl_csr_writedata_1;
input 	avl_csr_writedata_2;
input 	avl_csr_writedata_3;
input 	avl_csr_writedata_4;
input 	avl_csr_writedata_5;
input 	avl_csr_writedata_6;
input 	avl_csr_writedata_7;
input 	avl_csr_writedata_8;
input 	avl_csr_writedata_9;
input 	avl_csr_writedata_10;
input 	avl_csr_writedata_11;
input 	avl_csr_writedata_12;
input 	avl_csr_writedata_13;
input 	avl_csr_writedata_14;
input 	avl_csr_writedata_15;
input 	avl_csr_writedata_16;
input 	avl_csr_writedata_17;
input 	avl_csr_writedata_18;
input 	avl_csr_writedata_19;
input 	avl_csr_writedata_20;
input 	avl_csr_writedata_21;
input 	avl_csr_writedata_22;
input 	avl_csr_writedata_23;
input 	avl_csr_writedata_24;
input 	avl_csr_writedata_25;
input 	avl_csr_writedata_26;
input 	avl_csr_writedata_27;
input 	avl_csr_writedata_28;
input 	avl_csr_writedata_29;
input 	avl_csr_writedata_30;
input 	avl_csr_writedata_31;
input 	avl_mem_read;
input 	avl_mem_burstcount_0;
input 	avl_mem_burstcount_6;
input 	avl_mem_burstcount_2;
input 	avl_mem_burstcount_1;
input 	avl_mem_burstcount_5;
input 	avl_mem_burstcount_4;
input 	avl_mem_burstcount_3;
input 	avl_mem_write;
input 	avl_mem_byteenable_0;
input 	avl_mem_byteenable_1;
input 	avl_mem_byteenable_2;
input 	avl_mem_byteenable_3;
input 	reset_reset;
input 	avl_mem_writedata_30;
input 	avl_mem_writedata_29;
input 	avl_mem_writedata_28;
input 	avl_mem_writedata_27;
input 	avl_mem_writedata_11;
input 	avl_mem_writedata_18;
input 	avl_mem_writedata_19;
input 	avl_mem_writedata_21;
input 	avl_mem_writedata_20;
input 	avl_mem_writedata_22;
input 	avl_mem_writedata_23;
input 	avl_mem_writedata_24;
input 	avl_mem_writedata_25;
input 	avl_mem_writedata_26;
input 	avl_mem_writedata_10;
input 	avl_mem_writedata_8;
input 	dut_asmiblock;
input 	avl_mem_writedata_13;
input 	avl_mem_writedata_17;
input 	avl_mem_writedata_16;
input 	avl_mem_writedata_15;
input 	avl_mem_writedata_31;
input 	avl_mem_writedata_14;
input 	avl_mem_writedata_9;
input 	avl_mem_address_6;
input 	avl_mem_address_14;
input 	avl_mem_writedata_0;
input 	avl_mem_address_10;
input 	avl_mem_address_18;
input 	avl_mem_address_2;
input 	avl_mem_writedata_4;
input 	avl_mem_writedata_12;
input 	avl_mem_address_8;
input 	avl_mem_address_16;
input 	avl_mem_address_0;
input 	avl_mem_writedata_2;
input 	avl_mem_address_15;
input 	avl_mem_address_7;
input 	avl_mem_writedata_1;
input 	avl_mem_address_17;
input 	avl_mem_address_9;
input 	avl_mem_address_1;
input 	avl_mem_writedata_3;
input 	avl_mem_address_19;
input 	avl_mem_address_11;
input 	avl_mem_address_3;
input 	avl_mem_writedata_5;
input 	avl_mem_address_12;
input 	avl_mem_address_20;
input 	avl_mem_address_4;
input 	avl_mem_writedata_6;
input 	avl_mem_address_13;
input 	avl_mem_address_5;
input 	avl_mem_writedata_7;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \serial_flash_inf_cmd_gen_inst|data_num_lines[1]~q ;
wire \serial_flash_inf_cmd_gen_inst|data_num_lines[2]~q ;
wire \serial_flash_inf_cmd_gen_inst|addr_num_lines[2]~q ;
wire \serial_flash_inf_cmd_gen_inst|addr_num_lines[1]~q ;
wire \csr_controller|state.ST_IDLE~q ;
wire \xip_controller|hold_waitrequest~q ;
wire \csr_controller|csr_wr_inst_data[0]~q ;
wire \csr_controller|csr_rd_inst_data[0]~q ;
wire \csr_controller|csr_op_protocol_data[0]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[0]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[0]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[0]~q ;
wire \csr_controller|csr_delay_setting_data[0]~q ;
wire \csr_controller|csr_clk_baud_rate_data[0]~q ;
wire \csr_controller|csr_control_data[0]~q ;
wire \csr_controller|csr_rd_capturing_data[0]~q ;
wire \rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \csr_controller|csr_wr_inst_data[1]~q ;
wire \csr_controller|csr_rd_inst_data[1]~q ;
wire \csr_controller|csr_op_protocol_data[1]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[1]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[1]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[1]~q ;
wire \csr_controller|csr_delay_setting_data[1]~q ;
wire \csr_controller|csr_clk_baud_rate_data[1]~q ;
wire \csr_controller|csr_rd_capturing_data[1]~q ;
wire \csr_controller|csr_wr_inst_data[2]~q ;
wire \csr_controller|csr_rd_inst_data[2]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[2]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[2]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[2]~q ;
wire \csr_controller|csr_delay_setting_data[2]~q ;
wire \csr_controller|csr_clk_baud_rate_data[2]~q ;
wire \csr_controller|csr_rd_capturing_data[2]~q ;
wire \csr_controller|csr_wr_inst_data[3]~q ;
wire \csr_controller|csr_rd_inst_data[3]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[3]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[3]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[3]~q ;
wire \csr_controller|csr_delay_setting_data[3]~q ;
wire \csr_controller|csr_clk_baud_rate_data[3]~q ;
wire \csr_controller|csr_rd_capturing_data[3]~q ;
wire \csr_controller|csr_wr_inst_data[4]~q ;
wire \csr_controller|csr_delay_setting_data[4]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[4]~q ;
wire \csr_controller|csr_op_protocol_data[4]~q ;
wire \csr_controller|csr_clk_baud_rate_data[4]~q ;
wire \csr_controller|csr_control_data[4]~q ;
wire \csr_controller|csr_rd_inst_data[4]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[4]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[4]~q ;
wire \csr_controller|csr_delay_setting_data[5]~q ;
wire \csr_controller|csr_wr_inst_data[5]~q ;
wire \csr_controller|csr_rd_inst_data[5]~q ;
wire \csr_controller|csr_op_protocol_data[5]~q ;
wire \csr_controller|csr_control_data[5]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[5]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[5]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[5]~q ;
wire \csr_controller|csr_wr_inst_data[6]~q ;
wire \csr_controller|csr_rd_inst_data[6]~q ;
wire \csr_controller|csr_delay_setting_data[6]~q ;
wire \csr_controller|csr_control_data[6]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[6]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[6]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[6]~q ;
wire \csr_controller|csr_delay_setting_data[7]~q ;
wire \csr_controller|csr_wr_inst_data[7]~q ;
wire \csr_controller|csr_rd_inst_data[7]~q ;
wire \csr_controller|csr_control_data[7]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[7]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[7]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[7]~q ;
wire \csr_controller|csr_rd_inst_data[8]~q ;
wire \csr_controller|csr_op_protocol_data[8]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[8]~q ;
wire \csr_controller|csr_control_data[8]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[8]~q ;
wire \csr_controller|csr_wr_inst_data[8]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[8]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[9]~q ;
wire \csr_controller|csr_rd_inst_data[9]~q ;
wire \csr_controller|csr_op_protocol_data[9]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[9]~q ;
wire \csr_controller|csr_wr_inst_data[9]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[9]~q ;
wire \csr_controller|csr_rd_inst_data[10]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[10]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[10]~q ;
wire \csr_controller|csr_wr_inst_data[10]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[10]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[11]~q ;
wire \csr_controller|csr_rd_inst_data[11]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[11]~q ;
wire \csr_controller|csr_wr_inst_data[11]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[11]~q ;
wire \csr_controller|csr_rd_inst_data[12]~q ;
wire \csr_controller|csr_op_protocol_data[12]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[12]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[12]~q ;
wire \csr_controller|csr_wr_inst_data[12]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[12]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[13]~q ;
wire \csr_controller|csr_op_protocol_data[13]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[13]~q ;
wire \csr_controller|csr_wr_inst_data[13]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[13]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[14]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[14]~q ;
wire \csr_controller|csr_wr_inst_data[14]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[14]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[15]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[15]~q ;
wire \csr_controller|csr_wr_inst_data[15]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[15]~q ;
wire \csr_controller|csr_op_protocol_data[16]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[16]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[16]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[16]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[17]~q ;
wire \csr_controller|csr_op_protocol_data[17]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[17]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[17]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[18]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[18]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[18]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[19]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[19]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[19]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[20]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[20]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[20]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[21]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[21]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[21]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[22]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[22]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[22]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[23]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[23]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[23]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[24]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[24]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[24]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[25]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[25]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[25]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[26]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[26]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[26]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[27]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[27]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[27]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[28]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[28]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[28]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[29]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[29]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[29]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[30]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[30]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[30]~q ;
wire \csr_controller|csr_flash_cmd_addr_data[31]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_0_data[31]~q ;
wire \csr_controller|csr_flash_cmd_wr_data_1_data[31]~q ;
wire \serial_flash_inf_cmd_gen_inst|state.ST_SEND_DUMMY_RSP~q ;
wire \serial_flash_inf_cmd_gen_inst|data_adapter_8_32_inst|out_valid~q ;
wire \serial_flash_inf_cmd_gen_inst|data_adapter_8_32_inst|out_endofpacket~q ;
wire \serial_flash_inf_cmd_gen_inst|in_cmd_channel_reg[1]~q ;
wire \csr_controller|state.ST_WAIT_RSP~q ;
wire \merlin_demultiplexer_0|sink_ready~0_combout ;
wire \serial_flash_inf_cmd_gen_inst|data_adapter_8_32_inst|out_data[0]~q ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[0]~0_combout ;
wire \xip_controller|current_state.STATE_READ_DATA~q ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[1]~1_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[2]~2_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[3]~3_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[4]~4_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[5]~5_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[6]~6_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[7]~7_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[8]~8_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[9]~9_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[10]~10_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[11]~11_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[12]~12_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[13]~13_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[14]~14_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[15]~15_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[16]~16_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[17]~17_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[18]~18_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[19]~19_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[20]~20_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[21]~21_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[22]~22_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[23]~23_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[24]~24_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[25]~25_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[26]~26_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[27]~27_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[28]~28_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[29]~29_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[30]~30_combout ;
wire \serial_flash_inf_cmd_gen_inst|out_rsp_data[31]~31_combout ;
wire \serial_flash_inf_cmd_gen_inst|in_cmd_channel_reg[0]~q ;
wire \serial_flash_inf_cmd_gen_inst|header_information[30]~q ;
wire \serial_flash_inf_cmd_gen_inst|header_information[29]~q ;
wire \serial_flash_inf_cmd_gen_inst|header_information[28]~q ;
wire \serial_flash_inf_cmd_gen_inst|header_information[27]~q ;
wire \merlin_demultiplexer_0|WideOr0~combout ;
wire \serial_flash_inf_cmd_gen_inst|state.ST_IDLE~q ;
wire \multiplexer|saved_grant[1]~q ;
wire \csr_controller|state.ST_SEND_HEADER~q ;
wire \multiplexer|saved_grant[0]~q ;
wire \xip_controller|current_state.STATE_WR_CMD~q ;
wire \xip_controller|current_state.STATE_STATUS_CMD~q ;
wire \xip_controller|current_state.STATE_POLL_CMD~q ;
wire \xip_controller|current_state.STATE_READ_CMD~q ;
wire \xip_controller|WideOr13~0_combout ;
wire \multiplexer|src_startofpacket~combout ;
wire \multiplexer|src_valid~0_combout ;
wire \xip_controller|current_state.STATE_WR_DATA~q ;
wire \xip_controller|cmd_valid~0_combout ;
wire \serial_flash_inf_cmd_gen_inst|state.ST_SEND_DATA~q ;
wire \serial_flash_inf_cmd_gen_inst|state.ST_SEND_ADDR~q ;
wire \serial_flash_inf_cmd_gen_inst|Selector18~2_combout ;
wire \serial_flash_inf_cmd_gen_inst|op_num_lines[1]~q ;
wire \serial_flash_inf_cmd_gen_inst|data_num_lines[0]~q ;
wire \serial_flash_inf_cmd_gen_inst|op_num_lines[0]~q ;
wire \qspi_inf_inst|demultiplexer_inst|WideOr0~3_combout ;
wire \qspi_inf_inst|adapter_8_4_inst|in_ready~combout ;
wire \serial_flash_inf_cmd_gen_inst|op_num_lines[2]~q ;
wire \qspi_inf_inst|demultiplexer_inst|WideOr0~4_combout ;
wire \serial_flash_inf_cmd_gen_inst|adap_out_cmd_ready~0_combout ;
wire \serial_flash_inf_cmd_gen_inst|Selector18~3_combout ;
wire \csr_controller|state.ST_SEND_DATA_1~q ;
wire \csr_controller|state.ST_SEND_DATA_0~q ;
wire \csr_controller|has_data_in~q ;
wire \csr_controller|more_than_4bytes_data~q ;
wire \multiplexer|src_payload[0]~1_combout ;
wire \serial_flash_inf_cmd_gen_inst|Selector18~5_combout ;
wire \multiplexer|sink0_ready~1_combout ;
wire \serial_flash_inf_cmd_gen_inst|header_information[11]~q ;
wire \multiplexer|src_data[30]~3_combout ;
wire \xip_controller|is_burst_reg~q ;
wire \xip_controller|mem_write_data_reg[30]~q ;
wire \xip_controller|mem_byteenable_reg[0]~q ;
wire \xip_controller|mem_byteenable_reg[3]~q ;
wire \xip_controller|mem_byteenable_reg[2]~q ;
wire \xip_controller|mem_byteenable_reg[1]~q ;
wire \multiplexer|src_data[30]~5_combout ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[30]~q ;
wire \xip_controller|cmd_valid~1_combout ;
wire \multiplexer|src_data[30]~7_combout ;
wire \multiplexer|src_data[30]~8_combout ;
wire \multiplexer|src_data[29]~10_combout ;
wire \xip_controller|mem_write_data_reg[29]~q ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[29]~q ;
wire \multiplexer|src_data[29]~12_combout ;
wire \multiplexer|src_data[29]~13_combout ;
wire \multiplexer|src_data[28]~15_combout ;
wire \xip_controller|mem_write_data_reg[28]~q ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[28]~q ;
wire \multiplexer|src_data[28]~17_combout ;
wire \multiplexer|src_data[28]~18_combout ;
wire \multiplexer|src_data[27]~20_combout ;
wire \xip_controller|mem_write_data_reg[27]~q ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[27]~q ;
wire \multiplexer|src_data[27]~22_combout ;
wire \multiplexer|src_data[27]~23_combout ;
wire \serial_flash_inf_cmd_gen_inst|state.ST_SEND_OPCODE~q ;
wire \serial_flash_inf_cmd_gen_inst|Selector8~0_combout ;
wire \qspi_inf_inst|demux_channel[2]~1_combout ;
wire \qspi_inf_inst|demultiplexer_inst|sink_ready~0_combout ;
wire \serial_flash_inf_cmd_gen_inst|addr_num_lines[0]~q ;
wire \qspi_inf_inst|demultiplexer_inst|WideOr0~5_combout ;
wire \qspi_inf_inst|out_rsp_valid~q ;
wire \multiplexer|WideOr1~combout ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[32]~q ;
wire \multiplexer|src_payload[0]~3_combout ;
wire \multiplexer|sink1_ready~combout ;
wire \qspi_inf_inst|demultiplexer_inst|WideOr0~7_combout ;
wire \qspi_inf_inst|demultiplexer_inst|WideOr0~8_combout ;
wire \qspi_inf_inst|demultiplexer_inst|WideOr0~11_combout ;
wire \csr_controller|Selector34~0_combout ;
wire \qspi_inf_inst|out_rsp_data[0]~q ;
wire \qspi_inf_inst|out_rsp_data[1]~q ;
wire \qspi_inf_inst|out_rsp_data[2]~q ;
wire \qspi_inf_inst|out_rsp_data[3]~q ;
wire \qspi_inf_inst|out_rsp_data[4]~q ;
wire \qspi_inf_inst|out_rsp_data[5]~q ;
wire \qspi_inf_inst|out_rsp_data[6]~q ;
wire \qspi_inf_inst|out_rsp_data[7]~q ;
wire \serial_flash_inf_cmd_gen_inst|header_information[13]~q ;
wire \serial_flash_inf_cmd_gen_inst|header_information[17]~q ;
wire \serial_flash_inf_cmd_gen_inst|header_information[16]~q ;
wire \serial_flash_inf_cmd_gen_inst|header_information[15]~q ;
wire \serial_flash_inf_cmd_gen_inst|header_information[14]~q ;
wire \csr_controller|has_data_out~q ;
wire \multiplexer|src_data[11]~25_combout ;
wire \xip_controller|cmd_data[11]~combout ;
wire \multiplexer|src_data[11]~26_combout ;
wire \csr_controller|numb_data[0]~q ;
wire \xip_controller|Add1~1_combout ;
wire \xip_controller|Selector20~0_combout ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[18]~q ;
wire \xip_controller|mem_write_data_reg[18]~q ;
wire \multiplexer|src_data[18]~32_combout ;
wire \csr_controller|numb_data[1]~q ;
wire \multiplexer|src_data[19]~34_combout ;
wire \xip_controller|Add1~2_combout ;
wire \xip_controller|mem_write_data_reg[19]~q ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[19]~q ;
wire \multiplexer|src_data[19]~37_combout ;
wire \multiplexer|src_data[19]~38_combout ;
wire \csr_controller|numb_data[3]~q ;
wire \multiplexer|src_data[21]~40_combout ;
wire \xip_controller|mem_write_data_reg[21]~q ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[21]~q ;
wire \xip_controller|mem_burstcount_reg[1]~q ;
wire \multiplexer|src_data[21]~43_combout ;
wire \multiplexer|src_data[21]~44_combout ;
wire \csr_controller|numb_data[2]~q ;
wire \multiplexer|src_data[20]~46_combout ;
wire \xip_controller|mem_write_data_reg[20]~q ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[20]~q ;
wire \xip_controller|mem_burstcount_reg[0]~q ;
wire \multiplexer|src_data[20]~50_combout ;
wire \multiplexer|src_data[20]~51_combout ;
wire \xip_controller|mem_write_data_reg[22]~q ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[22]~q ;
wire \xip_controller|mem_burstcount_reg[2]~q ;
wire \multiplexer|src_data[22]~55_combout ;
wire \xip_controller|mem_write_data_reg[23]~q ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[23]~q ;
wire \xip_controller|mem_burstcount_reg[3]~q ;
wire \multiplexer|src_data[23]~59_combout ;
wire \xip_controller|mem_write_data_reg[24]~q ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[24]~q ;
wire \xip_controller|mem_burstcount_reg[4]~q ;
wire \multiplexer|src_data[24]~63_combout ;
wire \xip_controller|mem_write_data_reg[25]~q ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[25]~q ;
wire \xip_controller|mem_burstcount_reg[5]~q ;
wire \multiplexer|src_data[25]~67_combout ;
wire \xip_controller|mem_write_data_reg[26]~q ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[26]~q ;
wire \xip_controller|mem_burstcount_reg[6]~q ;
wire \multiplexer|src_data[26]~71_combout ;
wire \qspi_inf_inst|demultiplexer_inst|WideOr0~13_combout ;
wire \multiplexer|src_data[10]~73_combout ;
wire \xip_controller|cmd_data[10]~combout ;
wire \multiplexer|src_data[10]~74_combout ;
wire \csr_controller|has_addr~q ;
wire \multiplexer|src_data[8]~76_combout ;
wire \xip_controller|cmd_data[8]~combout ;
wire \multiplexer|src_data[8]~77_combout ;
wire \csr_controller|numb_dummy[0]~q ;
wire \multiplexer|src_data[13]~79_combout ;
wire \xip_controller|cmd_data[13]~combout ;
wire \multiplexer|src_data[13]~80_combout ;
wire \csr_controller|numb_dummy[4]~q ;
wire \multiplexer|src_data[17]~82_combout ;
wire \xip_controller|mem_write_data_reg[17]~q ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[17]~q ;
wire \multiplexer|src_data[17]~84_combout ;
wire \multiplexer|src_data[17]~85_combout ;
wire \csr_controller|numb_dummy[3]~q ;
wire \multiplexer|src_data[16]~87_combout ;
wire \xip_controller|mem_write_data_reg[16]~q ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[16]~q ;
wire \multiplexer|src_data[16]~89_combout ;
wire \multiplexer|src_data[16]~90_combout ;
wire \csr_controller|numb_dummy[2]~q ;
wire \multiplexer|src_data[15]~92_combout ;
wire \xip_controller|mem_write_data_reg[31]~q ;
wire \xip_controller|cmd_data[15]~combout ;
wire \multiplexer|src_data[15]~93_combout ;
wire \csr_controller|numb_dummy[1]~q ;
wire \multiplexer|src_data[14]~95_combout ;
wire \xip_controller|cmd_data[14]~combout ;
wire \multiplexer|src_data[14]~96_combout ;
wire \csr_controller|is_4bytes_addr~q ;
wire \multiplexer|src_data[9]~98_combout ;
wire \xip_controller|cmd_data[9]~combout ;
wire \multiplexer|src_data[9]~99_combout ;
wire \serial_flash_inf_cmd_gen_inst|Selector20~2_combout ;
wire \serial_flash_inf_cmd_gen_inst|Selector16~3_combout ;
wire \serial_flash_inf_cmd_gen_inst|Selector12~3_combout ;
wire \serial_flash_inf_cmd_gen_inst|Selector14~3_combout ;
wire \serial_flash_inf_cmd_gen_inst|Selector15~3_combout ;
wire \serial_flash_inf_cmd_gen_inst|Selector13~3_combout ;
wire \serial_flash_inf_cmd_gen_inst|Selector11~3_combout ;
wire \serial_flash_inf_cmd_gen_inst|Selector10~3_combout ;
wire \serial_flash_inf_cmd_gen_inst|Selector9~4_combout ;
wire \serial_flash_inf_cmd_gen_inst|Selector17~0_combout ;
wire \xip_controller|mem_addr_reg[6]~q ;
wire \xip_controller|mem_addr_reg[14]~q ;
wire \xip_controller|addr_bytes_xip[0]~0_combout ;
wire \csr_controller|opcode[0]~q ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[0]~q ;
wire \xip_controller|cmd_data[0]~36_combout ;
wire \multiplexer|src_data[0]~102_combout ;
wire \xip_controller|mem_addr_reg[10]~q ;
wire \xip_controller|mem_addr_reg[18]~q ;
wire \xip_controller|mem_addr_reg[2]~q ;
wire \csr_controller|opcode[4]~q ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[4]~q ;
wire \xip_controller|cmd_data[4]~43_combout ;
wire \multiplexer|src_data[4]~105_combout ;
wire \xip_controller|mem_addr_reg[8]~q ;
wire \xip_controller|mem_addr_reg[16]~q ;
wire \xip_controller|mem_addr_reg[0]~q ;
wire \csr_controller|opcode[2]~q ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[2]~q ;
wire \xip_controller|cmd_data[2]~50_combout ;
wire \multiplexer|src_data[2]~108_combout ;
wire \xip_controller|mem_addr_reg[15]~q ;
wire \xip_controller|mem_addr_reg[7]~q ;
wire \xip_controller|WideOr19~0_combout ;
wire \csr_controller|opcode[1]~q ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[1]~q ;
wire \xip_controller|cmd_data[1]~57_combout ;
wire \multiplexer|src_data[1]~111_combout ;
wire \xip_controller|mem_addr_reg[17]~q ;
wire \xip_controller|mem_addr_reg[9]~q ;
wire \xip_controller|mem_addr_reg[1]~q ;
wire \csr_controller|opcode[3]~q ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[3]~q ;
wire \xip_controller|cmd_data[3]~64_combout ;
wire \multiplexer|src_data[3]~114_combout ;
wire \xip_controller|mem_addr_reg[19]~q ;
wire \xip_controller|mem_addr_reg[11]~q ;
wire \xip_controller|mem_addr_reg[3]~q ;
wire \csr_controller|opcode[5]~q ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[5]~q ;
wire \xip_controller|cmd_data[5]~71_combout ;
wire \multiplexer|src_data[5]~117_combout ;
wire \xip_controller|mem_addr_reg[12]~q ;
wire \xip_controller|mem_addr_reg[20]~q ;
wire \xip_controller|mem_addr_reg[4]~q ;
wire \csr_controller|opcode[6]~q ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[6]~q ;
wire \xip_controller|cmd_data[6]~78_combout ;
wire \multiplexer|src_data[6]~120_combout ;
wire \xip_controller|mem_addr_reg[13]~q ;
wire \xip_controller|mem_addr_reg[5]~q ;
wire \csr_controller|opcode[7]~q ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[7]~q ;
wire \xip_controller|cmd_data[7]~85_combout ;
wire \multiplexer|src_data[7]~123_combout ;
wire \csr_controller|has_dummy~q ;
wire \xip_controller|cmd_data[12]~combout ;
wire \xip_controller|avst_fifo_inst|avst_fifo|out_payload[31]~q ;


flashLoader_altera_reset_controller rst_controller(
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk_clk(clk_clk),
	.reset_reset(reset_reset));

flashLoader_flashLoader_intel_generic_serial_flash_interface_top_0_qspi_inf_inst qspi_inf_inst(
	.data_num_lines_1(\serial_flash_inf_cmd_gen_inst|data_num_lines[1]~q ),
	.data_num_lines_2(\serial_flash_inf_cmd_gen_inst|data_num_lines[2]~q ),
	.addr_num_lines_2(\serial_flash_inf_cmd_gen_inst|addr_num_lines[2]~q ),
	.addr_num_lines_1(\serial_flash_inf_cmd_gen_inst|addr_num_lines[1]~q ),
	.flash_clk_reg1(flash_clk_reg),
	.oe_reg1(oe_reg),
	.ncs_reg_0(ncs_reg_0),
	.flash_data_out_reg_0(flash_data_out_reg_0),
	.csr_delay_setting_data_0(\csr_controller|csr_delay_setting_data[0]~q ),
	.csr_clk_baud_rate_data_0(\csr_controller|csr_clk_baud_rate_data[0]~q ),
	.qspi_interface_en(\csr_controller|csr_control_data[0]~q ),
	.csr_rd_capturing_data_0(\csr_controller|csr_rd_capturing_data[0]~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.csr_delay_setting_data_1(\csr_controller|csr_delay_setting_data[1]~q ),
	.csr_clk_baud_rate_data_1(\csr_controller|csr_clk_baud_rate_data[1]~q ),
	.csr_rd_capturing_data_1(\csr_controller|csr_rd_capturing_data[1]~q ),
	.csr_delay_setting_data_2(\csr_controller|csr_delay_setting_data[2]~q ),
	.csr_clk_baud_rate_data_2(\csr_controller|csr_clk_baud_rate_data[2]~q ),
	.csr_rd_capturing_data_2(\csr_controller|csr_rd_capturing_data[2]~q ),
	.csr_delay_setting_data_3(\csr_controller|csr_delay_setting_data[3]~q ),
	.csr_clk_baud_rate_data_3(\csr_controller|csr_clk_baud_rate_data[3]~q ),
	.csr_rd_capturing_data_3(\csr_controller|csr_rd_capturing_data[3]~q ),
	.csr_delay_setting_data_4(\csr_controller|csr_delay_setting_data[4]~q ),
	.csr_clk_baud_rate_data_4(\csr_controller|csr_clk_baud_rate_data[4]~q ),
	.csr_delay_setting_data_5(\csr_controller|csr_delay_setting_data[5]~q ),
	.csr_delay_setting_data_6(\csr_controller|csr_delay_setting_data[6]~q ),
	.csr_delay_setting_data_7(\csr_controller|csr_delay_setting_data[7]~q ),
	.in_cmd_channel_reg_1(\serial_flash_inf_cmd_gen_inst|in_cmd_channel_reg[1]~q ),
	.in_cmd_channel_reg_0(\serial_flash_inf_cmd_gen_inst|in_cmd_channel_reg[0]~q ),
	.header_information_30(\serial_flash_inf_cmd_gen_inst|header_information[30]~q ),
	.header_information_29(\serial_flash_inf_cmd_gen_inst|header_information[29]~q ),
	.header_information_28(\serial_flash_inf_cmd_gen_inst|header_information[28]~q ),
	.header_information_27(\serial_flash_inf_cmd_gen_inst|header_information[27]~q ),
	.stateST_IDLE(\serial_flash_inf_cmd_gen_inst|state.ST_IDLE~q ),
	.stateST_SEND_DATA(\serial_flash_inf_cmd_gen_inst|state.ST_SEND_DATA~q ),
	.stateST_SEND_ADDR(\serial_flash_inf_cmd_gen_inst|state.ST_SEND_ADDR~q ),
	.op_num_lines_1(\serial_flash_inf_cmd_gen_inst|op_num_lines[1]~q ),
	.data_num_lines_0(\serial_flash_inf_cmd_gen_inst|data_num_lines[0]~q ),
	.op_num_lines_0(\serial_flash_inf_cmd_gen_inst|op_num_lines[0]~q ),
	.WideOr0(\qspi_inf_inst|demultiplexer_inst|WideOr0~3_combout ),
	.in_ready(\qspi_inf_inst|adapter_8_4_inst|in_ready~combout ),
	.op_num_lines_2(\serial_flash_inf_cmd_gen_inst|op_num_lines[2]~q ),
	.WideOr01(\qspi_inf_inst|demultiplexer_inst|WideOr0~4_combout ),
	.header_information_11(\serial_flash_inf_cmd_gen_inst|header_information[11]~q ),
	.stateST_SEND_OPCODE(\serial_flash_inf_cmd_gen_inst|state.ST_SEND_OPCODE~q ),
	.Selector8(\serial_flash_inf_cmd_gen_inst|Selector8~0_combout ),
	.demux_channel_2(\qspi_inf_inst|demux_channel[2]~1_combout ),
	.in_cmd_ready(\qspi_inf_inst|demultiplexer_inst|sink_ready~0_combout ),
	.addr_num_lines_0(\serial_flash_inf_cmd_gen_inst|addr_num_lines[0]~q ),
	.WideOr02(\qspi_inf_inst|demultiplexer_inst|WideOr0~5_combout ),
	.out_rsp_valid1(\qspi_inf_inst|out_rsp_valid~q ),
	.WideOr03(\qspi_inf_inst|demultiplexer_inst|WideOr0~7_combout ),
	.WideOr04(\qspi_inf_inst|demultiplexer_inst|WideOr0~8_combout ),
	.WideOr05(\qspi_inf_inst|demultiplexer_inst|WideOr0~11_combout ),
	.out_rsp_data_0(\qspi_inf_inst|out_rsp_data[0]~q ),
	.out_rsp_data_1(\qspi_inf_inst|out_rsp_data[1]~q ),
	.out_rsp_data_2(\qspi_inf_inst|out_rsp_data[2]~q ),
	.out_rsp_data_3(\qspi_inf_inst|out_rsp_data[3]~q ),
	.out_rsp_data_4(\qspi_inf_inst|out_rsp_data[4]~q ),
	.out_rsp_data_5(\qspi_inf_inst|out_rsp_data[5]~q ),
	.out_rsp_data_6(\qspi_inf_inst|out_rsp_data[6]~q ),
	.out_rsp_data_7(\qspi_inf_inst|out_rsp_data[7]~q ),
	.header_information_13(\serial_flash_inf_cmd_gen_inst|header_information[13]~q ),
	.header_information_17(\serial_flash_inf_cmd_gen_inst|header_information[17]~q ),
	.header_information_16(\serial_flash_inf_cmd_gen_inst|header_information[16]~q ),
	.header_information_15(\serial_flash_inf_cmd_gen_inst|header_information[15]~q ),
	.header_information_14(\serial_flash_inf_cmd_gen_inst|header_information[14]~q ),
	.WideOr06(\qspi_inf_inst|demultiplexer_inst|WideOr0~13_combout ),
	.Selector20(\serial_flash_inf_cmd_gen_inst|Selector20~2_combout ),
	.Selector16(\serial_flash_inf_cmd_gen_inst|Selector16~3_combout ),
	.Selector12(\serial_flash_inf_cmd_gen_inst|Selector12~3_combout ),
	.Selector14(\serial_flash_inf_cmd_gen_inst|Selector14~3_combout ),
	.Selector15(\serial_flash_inf_cmd_gen_inst|Selector15~3_combout ),
	.Selector13(\serial_flash_inf_cmd_gen_inst|Selector13~3_combout ),
	.Selector11(\serial_flash_inf_cmd_gen_inst|Selector11~3_combout ),
	.Selector10(\serial_flash_inf_cmd_gen_inst|Selector10~3_combout ),
	.Selector9(\serial_flash_inf_cmd_gen_inst|Selector9~4_combout ),
	.Selector17(\serial_flash_inf_cmd_gen_inst|Selector17~0_combout ),
	.clk_clk(clk_clk),
	.dut_asmiblock(dut_asmiblock));

flashLoader_intel_generic_serial_flash_interface_cmd serial_flash_inf_cmd_gen_inst(
	.data_num_lines_1(\serial_flash_inf_cmd_gen_inst|data_num_lines[1]~q ),
	.data_num_lines_2(\serial_flash_inf_cmd_gen_inst|data_num_lines[2]~q ),
	.addr_num_lines_2(\serial_flash_inf_cmd_gen_inst|addr_num_lines[2]~q ),
	.addr_num_lines_1(\serial_flash_inf_cmd_gen_inst|addr_num_lines[1]~q ),
	.csr_op_protocol_data_0(\csr_controller|csr_op_protocol_data[0]~q ),
	.csr_flash_cmd_addr_data_0(\csr_controller|csr_flash_cmd_addr_data[0]~q ),
	.reset(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.csr_op_protocol_data_1(\csr_controller|csr_op_protocol_data[1]~q ),
	.csr_flash_cmd_addr_data_1(\csr_controller|csr_flash_cmd_addr_data[1]~q ),
	.csr_flash_cmd_addr_data_2(\csr_controller|csr_flash_cmd_addr_data[2]~q ),
	.csr_flash_cmd_addr_data_3(\csr_controller|csr_flash_cmd_addr_data[3]~q ),
	.csr_flash_cmd_addr_data_4(\csr_controller|csr_flash_cmd_addr_data[4]~q ),
	.csr_op_protocol_data_4(\csr_controller|csr_op_protocol_data[4]~q ),
	.csr_op_protocol_data_5(\csr_controller|csr_op_protocol_data[5]~q ),
	.csr_flash_cmd_addr_data_5(\csr_controller|csr_flash_cmd_addr_data[5]~q ),
	.csr_flash_cmd_addr_data_6(\csr_controller|csr_flash_cmd_addr_data[6]~q ),
	.csr_flash_cmd_addr_data_7(\csr_controller|csr_flash_cmd_addr_data[7]~q ),
	.csr_op_protocol_data_8(\csr_controller|csr_op_protocol_data[8]~q ),
	.csr_flash_cmd_addr_data_8(\csr_controller|csr_flash_cmd_addr_data[8]~q ),
	.csr_flash_cmd_addr_data_9(\csr_controller|csr_flash_cmd_addr_data[9]~q ),
	.csr_op_protocol_data_9(\csr_controller|csr_op_protocol_data[9]~q ),
	.csr_flash_cmd_addr_data_10(\csr_controller|csr_flash_cmd_addr_data[10]~q ),
	.csr_flash_cmd_addr_data_11(\csr_controller|csr_flash_cmd_addr_data[11]~q ),
	.csr_op_protocol_data_12(\csr_controller|csr_op_protocol_data[12]~q ),
	.csr_flash_cmd_addr_data_12(\csr_controller|csr_flash_cmd_addr_data[12]~q ),
	.csr_flash_cmd_wr_data_0_data_12(\csr_controller|csr_flash_cmd_wr_data_0_data[12]~q ),
	.csr_flash_cmd_wr_data_1_data_12(\csr_controller|csr_flash_cmd_wr_data_1_data[12]~q ),
	.csr_flash_cmd_addr_data_13(\csr_controller|csr_flash_cmd_addr_data[13]~q ),
	.csr_op_protocol_data_13(\csr_controller|csr_op_protocol_data[13]~q ),
	.csr_flash_cmd_addr_data_14(\csr_controller|csr_flash_cmd_addr_data[14]~q ),
	.csr_flash_cmd_addr_data_15(\csr_controller|csr_flash_cmd_addr_data[15]~q ),
	.csr_op_protocol_data_16(\csr_controller|csr_op_protocol_data[16]~q ),
	.csr_flash_cmd_addr_data_16(\csr_controller|csr_flash_cmd_addr_data[16]~q ),
	.csr_flash_cmd_addr_data_17(\csr_controller|csr_flash_cmd_addr_data[17]~q ),
	.csr_op_protocol_data_17(\csr_controller|csr_op_protocol_data[17]~q ),
	.csr_flash_cmd_addr_data_18(\csr_controller|csr_flash_cmd_addr_data[18]~q ),
	.csr_flash_cmd_addr_data_19(\csr_controller|csr_flash_cmd_addr_data[19]~q ),
	.csr_flash_cmd_addr_data_20(\csr_controller|csr_flash_cmd_addr_data[20]~q ),
	.csr_flash_cmd_addr_data_21(\csr_controller|csr_flash_cmd_addr_data[21]~q ),
	.csr_flash_cmd_addr_data_22(\csr_controller|csr_flash_cmd_addr_data[22]~q ),
	.csr_flash_cmd_addr_data_23(\csr_controller|csr_flash_cmd_addr_data[23]~q ),
	.csr_flash_cmd_addr_data_24(\csr_controller|csr_flash_cmd_addr_data[24]~q ),
	.csr_flash_cmd_addr_data_25(\csr_controller|csr_flash_cmd_addr_data[25]~q ),
	.csr_flash_cmd_addr_data_26(\csr_controller|csr_flash_cmd_addr_data[26]~q ),
	.csr_flash_cmd_addr_data_27(\csr_controller|csr_flash_cmd_addr_data[27]~q ),
	.csr_flash_cmd_addr_data_28(\csr_controller|csr_flash_cmd_addr_data[28]~q ),
	.csr_flash_cmd_addr_data_29(\csr_controller|csr_flash_cmd_addr_data[29]~q ),
	.csr_flash_cmd_addr_data_30(\csr_controller|csr_flash_cmd_addr_data[30]~q ),
	.csr_flash_cmd_addr_data_31(\csr_controller|csr_flash_cmd_addr_data[31]~q ),
	.csr_flash_cmd_wr_data_0_data_31(\csr_controller|csr_flash_cmd_wr_data_0_data[31]~q ),
	.csr_flash_cmd_wr_data_1_data_31(\csr_controller|csr_flash_cmd_wr_data_1_data[31]~q ),
	.stateST_SEND_DUMMY_RSP(\serial_flash_inf_cmd_gen_inst|state.ST_SEND_DUMMY_RSP~q ),
	.out_valid(\serial_flash_inf_cmd_gen_inst|data_adapter_8_32_inst|out_valid~q ),
	.out_endofpacket(\serial_flash_inf_cmd_gen_inst|data_adapter_8_32_inst|out_endofpacket~q ),
	.in_cmd_channel_reg_1(\serial_flash_inf_cmd_gen_inst|in_cmd_channel_reg[1]~q ),
	.stateST_WAIT_RSP(\csr_controller|state.ST_WAIT_RSP~q ),
	.out_data_0(\serial_flash_inf_cmd_gen_inst|data_adapter_8_32_inst|out_data[0]~q ),
	.out_rsp_data_0(\serial_flash_inf_cmd_gen_inst|out_rsp_data[0]~0_combout ),
	.current_stateSTATE_READ_DATA(\xip_controller|current_state.STATE_READ_DATA~q ),
	.out_rsp_data_1(\serial_flash_inf_cmd_gen_inst|out_rsp_data[1]~1_combout ),
	.out_rsp_data_2(\serial_flash_inf_cmd_gen_inst|out_rsp_data[2]~2_combout ),
	.out_rsp_data_3(\serial_flash_inf_cmd_gen_inst|out_rsp_data[3]~3_combout ),
	.out_rsp_data_4(\serial_flash_inf_cmd_gen_inst|out_rsp_data[4]~4_combout ),
	.out_rsp_data_5(\serial_flash_inf_cmd_gen_inst|out_rsp_data[5]~5_combout ),
	.out_rsp_data_6(\serial_flash_inf_cmd_gen_inst|out_rsp_data[6]~6_combout ),
	.out_rsp_data_7(\serial_flash_inf_cmd_gen_inst|out_rsp_data[7]~7_combout ),
	.out_rsp_data_8(\serial_flash_inf_cmd_gen_inst|out_rsp_data[8]~8_combout ),
	.out_rsp_data_9(\serial_flash_inf_cmd_gen_inst|out_rsp_data[9]~9_combout ),
	.out_rsp_data_10(\serial_flash_inf_cmd_gen_inst|out_rsp_data[10]~10_combout ),
	.out_rsp_data_11(\serial_flash_inf_cmd_gen_inst|out_rsp_data[11]~11_combout ),
	.out_rsp_data_12(\serial_flash_inf_cmd_gen_inst|out_rsp_data[12]~12_combout ),
	.out_rsp_data_13(\serial_flash_inf_cmd_gen_inst|out_rsp_data[13]~13_combout ),
	.out_rsp_data_14(\serial_flash_inf_cmd_gen_inst|out_rsp_data[14]~14_combout ),
	.out_rsp_data_15(\serial_flash_inf_cmd_gen_inst|out_rsp_data[15]~15_combout ),
	.out_rsp_data_16(\serial_flash_inf_cmd_gen_inst|out_rsp_data[16]~16_combout ),
	.out_rsp_data_17(\serial_flash_inf_cmd_gen_inst|out_rsp_data[17]~17_combout ),
	.out_rsp_data_18(\serial_flash_inf_cmd_gen_inst|out_rsp_data[18]~18_combout ),
	.out_rsp_data_19(\serial_flash_inf_cmd_gen_inst|out_rsp_data[19]~19_combout ),
	.out_rsp_data_20(\serial_flash_inf_cmd_gen_inst|out_rsp_data[20]~20_combout ),
	.out_rsp_data_21(\serial_flash_inf_cmd_gen_inst|out_rsp_data[21]~21_combout ),
	.out_rsp_data_22(\serial_flash_inf_cmd_gen_inst|out_rsp_data[22]~22_combout ),
	.out_rsp_data_23(\serial_flash_inf_cmd_gen_inst|out_rsp_data[23]~23_combout ),
	.out_rsp_data_24(\serial_flash_inf_cmd_gen_inst|out_rsp_data[24]~24_combout ),
	.out_rsp_data_25(\serial_flash_inf_cmd_gen_inst|out_rsp_data[25]~25_combout ),
	.out_rsp_data_26(\serial_flash_inf_cmd_gen_inst|out_rsp_data[26]~26_combout ),
	.out_rsp_data_27(\serial_flash_inf_cmd_gen_inst|out_rsp_data[27]~27_combout ),
	.out_rsp_data_28(\serial_flash_inf_cmd_gen_inst|out_rsp_data[28]~28_combout ),
	.out_rsp_data_29(\serial_flash_inf_cmd_gen_inst|out_rsp_data[29]~29_combout ),
	.out_rsp_data_30(\serial_flash_inf_cmd_gen_inst|out_rsp_data[30]~30_combout ),
	.out_rsp_data_31(\serial_flash_inf_cmd_gen_inst|out_rsp_data[31]~31_combout ),
	.in_cmd_channel_reg_0(\serial_flash_inf_cmd_gen_inst|in_cmd_channel_reg[0]~q ),
	.header_information_30(\serial_flash_inf_cmd_gen_inst|header_information[30]~q ),
	.header_information_29(\serial_flash_inf_cmd_gen_inst|header_information[29]~q ),
	.header_information_28(\serial_flash_inf_cmd_gen_inst|header_information[28]~q ),
	.header_information_27(\serial_flash_inf_cmd_gen_inst|header_information[27]~q ),
	.WideOr0(\merlin_demultiplexer_0|WideOr0~combout ),
	.stateST_IDLE(\serial_flash_inf_cmd_gen_inst|state.ST_IDLE~q ),
	.in_cmd_channel({\multiplexer|saved_grant[1]~q ,\multiplexer|saved_grant[0]~q }),
	.stateST_SEND_HEADER(\csr_controller|state.ST_SEND_HEADER~q ),
	.current_stateSTATE_WR_CMD(\xip_controller|current_state.STATE_WR_CMD~q ),
	.current_stateSTATE_READ_CMD(\xip_controller|current_state.STATE_READ_CMD~q ),
	.src_startofpacket(\multiplexer|src_startofpacket~combout ),
	.src_valid(\multiplexer|src_valid~0_combout ),
	.current_stateSTATE_WR_DATA(\xip_controller|current_state.STATE_WR_DATA~q ),
	.cmd_valid(\xip_controller|cmd_valid~0_combout ),
	.stateST_SEND_DATA(\serial_flash_inf_cmd_gen_inst|state.ST_SEND_DATA~q ),
	.stateST_SEND_ADDR(\serial_flash_inf_cmd_gen_inst|state.ST_SEND_ADDR~q ),
	.Selector18(\serial_flash_inf_cmd_gen_inst|Selector18~2_combout ),
	.op_num_lines_1(\serial_flash_inf_cmd_gen_inst|op_num_lines[1]~q ),
	.data_num_lines_0(\serial_flash_inf_cmd_gen_inst|data_num_lines[0]~q ),
	.op_num_lines_0(\serial_flash_inf_cmd_gen_inst|op_num_lines[0]~q ),
	.WideOr01(\qspi_inf_inst|demultiplexer_inst|WideOr0~3_combout ),
	.in_ready(\qspi_inf_inst|adapter_8_4_inst|in_ready~combout ),
	.op_num_lines_2(\serial_flash_inf_cmd_gen_inst|op_num_lines[2]~q ),
	.WideOr02(\qspi_inf_inst|demultiplexer_inst|WideOr0~4_combout ),
	.adap_out_cmd_ready(\serial_flash_inf_cmd_gen_inst|adap_out_cmd_ready~0_combout ),
	.Selector181(\serial_flash_inf_cmd_gen_inst|Selector18~3_combout ),
	.stateST_SEND_DATA_1(\csr_controller|state.ST_SEND_DATA_1~q ),
	.stateST_SEND_DATA_0(\csr_controller|state.ST_SEND_DATA_0~q ),
	.Selector182(\serial_flash_inf_cmd_gen_inst|Selector18~5_combout ),
	.header_information_11(\serial_flash_inf_cmd_gen_inst|header_information[11]~q ),
	.src_data_30(\multiplexer|src_data[30]~3_combout ),
	.is_burst_reg(\xip_controller|is_burst_reg~q ),
	.src_data_301(\multiplexer|src_data[30]~5_combout ),
	.src_data_302(\multiplexer|src_data[30]~7_combout ),
	.in_cmd_data({gnd,\multiplexer|src_data[30]~8_combout ,\multiplexer|src_data[29]~13_combout ,\multiplexer|src_data[28]~18_combout ,\multiplexer|src_data[27]~23_combout ,\multiplexer|src_data[26]~71_combout ,\multiplexer|src_data[25]~67_combout ,
\multiplexer|src_data[24]~63_combout ,\multiplexer|src_data[23]~59_combout ,\multiplexer|src_data[22]~55_combout ,\multiplexer|src_data[21]~44_combout ,\multiplexer|src_data[20]~51_combout ,\multiplexer|src_data[19]~38_combout ,
\multiplexer|src_data[18]~32_combout ,\multiplexer|src_data[17]~85_combout ,\multiplexer|src_data[16]~90_combout ,\multiplexer|src_data[15]~93_combout ,\multiplexer|src_data[14]~96_combout ,\multiplexer|src_data[13]~80_combout ,gnd,
\multiplexer|src_data[11]~26_combout ,\multiplexer|src_data[10]~74_combout ,\multiplexer|src_data[9]~99_combout ,\multiplexer|src_data[8]~77_combout ,\multiplexer|src_data[7]~123_combout ,\multiplexer|src_data[6]~120_combout ,
\multiplexer|src_data[5]~117_combout ,\multiplexer|src_data[4]~105_combout ,\multiplexer|src_data[3]~114_combout ,\multiplexer|src_data[2]~108_combout ,\multiplexer|src_data[1]~111_combout ,\multiplexer|src_data[0]~102_combout }),
	.src_data_29(\multiplexer|src_data[29]~10_combout ),
	.src_data_291(\multiplexer|src_data[29]~12_combout ),
	.src_data_28(\multiplexer|src_data[28]~15_combout ),
	.src_data_281(\multiplexer|src_data[28]~17_combout ),
	.src_data_27(\multiplexer|src_data[27]~20_combout ),
	.src_data_271(\multiplexer|src_data[27]~22_combout ),
	.stateST_SEND_OPCODE(\serial_flash_inf_cmd_gen_inst|state.ST_SEND_OPCODE~q ),
	.Selector8(\serial_flash_inf_cmd_gen_inst|Selector8~0_combout ),
	.demux_channel_2(\qspi_inf_inst|demux_channel[2]~1_combout ),
	.sink_ready(\qspi_inf_inst|demultiplexer_inst|sink_ready~0_combout ),
	.addr_num_lines_0(\serial_flash_inf_cmd_gen_inst|addr_num_lines[0]~q ),
	.WideOr03(\qspi_inf_inst|demultiplexer_inst|WideOr0~5_combout ),
	.out_rsp_valid(\qspi_inf_inst|out_rsp_valid~q ),
	.WideOr1(\multiplexer|WideOr1~combout ),
	.src_payload_0(\multiplexer|src_payload[0]~3_combout ),
	.WideOr04(\qspi_inf_inst|demultiplexer_inst|WideOr0~7_combout ),
	.WideOr05(\qspi_inf_inst|demultiplexer_inst|WideOr0~8_combout ),
	.WideOr06(\qspi_inf_inst|demultiplexer_inst|WideOr0~11_combout ),
	.out_rsp_data_01(\qspi_inf_inst|out_rsp_data[0]~q ),
	.out_rsp_data_110(\qspi_inf_inst|out_rsp_data[1]~q ),
	.out_rsp_data_210(\qspi_inf_inst|out_rsp_data[2]~q ),
	.out_rsp_data_32(\qspi_inf_inst|out_rsp_data[3]~q ),
	.out_rsp_data_41(\qspi_inf_inst|out_rsp_data[4]~q ),
	.out_rsp_data_51(\qspi_inf_inst|out_rsp_data[5]~q ),
	.out_rsp_data_61(\qspi_inf_inst|out_rsp_data[6]~q ),
	.out_rsp_data_71(\qspi_inf_inst|out_rsp_data[7]~q ),
	.header_information_13(\serial_flash_inf_cmd_gen_inst|header_information[13]~q ),
	.header_information_17(\serial_flash_inf_cmd_gen_inst|header_information[17]~q ),
	.header_information_16(\serial_flash_inf_cmd_gen_inst|header_information[16]~q ),
	.header_information_15(\serial_flash_inf_cmd_gen_inst|header_information[15]~q ),
	.header_information_14(\serial_flash_inf_cmd_gen_inst|header_information[14]~q ),
	.src_data_11(\multiplexer|src_data[11]~25_combout ),
	.cmd_data_11(\xip_controller|cmd_data[11]~combout ),
	.src_data_19(\multiplexer|src_data[19]~34_combout ),
	.src_data_191(\multiplexer|src_data[19]~37_combout ),
	.src_data_21(\multiplexer|src_data[21]~40_combout ),
	.src_data_211(\multiplexer|src_data[21]~43_combout ),
	.src_data_20(\multiplexer|src_data[20]~46_combout ),
	.src_data_201(\multiplexer|src_data[20]~50_combout ),
	.WideOr07(\qspi_inf_inst|demultiplexer_inst|WideOr0~13_combout ),
	.src_data_10(\multiplexer|src_data[10]~73_combout ),
	.cmd_data_10(\xip_controller|cmd_data[10]~combout ),
	.has_addr(\csr_controller|has_addr~q ),
	.src_data_8(\multiplexer|src_data[8]~76_combout ),
	.cmd_data_8(\xip_controller|cmd_data[8]~combout ),
	.src_data_13(\multiplexer|src_data[13]~79_combout ),
	.cmd_data_13(\xip_controller|cmd_data[13]~combout ),
	.src_data_17(\multiplexer|src_data[17]~82_combout ),
	.src_data_171(\multiplexer|src_data[17]~84_combout ),
	.src_data_16(\multiplexer|src_data[16]~87_combout ),
	.src_data_161(\multiplexer|src_data[16]~89_combout ),
	.src_data_15(\multiplexer|src_data[15]~92_combout ),
	.mem_write_data_reg_31(\xip_controller|mem_write_data_reg[31]~q ),
	.cmd_data_15(\xip_controller|cmd_data[15]~combout ),
	.src_data_14(\multiplexer|src_data[14]~95_combout ),
	.cmd_data_14(\xip_controller|cmd_data[14]~combout ),
	.src_data_9(\multiplexer|src_data[9]~98_combout ),
	.cmd_data_9(\xip_controller|cmd_data[9]~combout ),
	.Selector20(\serial_flash_inf_cmd_gen_inst|Selector20~2_combout ),
	.Selector16(\serial_flash_inf_cmd_gen_inst|Selector16~3_combout ),
	.Selector12(\serial_flash_inf_cmd_gen_inst|Selector12~3_combout ),
	.Selector14(\serial_flash_inf_cmd_gen_inst|Selector14~3_combout ),
	.Selector15(\serial_flash_inf_cmd_gen_inst|Selector15~3_combout ),
	.Selector13(\serial_flash_inf_cmd_gen_inst|Selector13~3_combout ),
	.Selector11(\serial_flash_inf_cmd_gen_inst|Selector11~3_combout ),
	.Selector10(\serial_flash_inf_cmd_gen_inst|Selector10~3_combout ),
	.Selector9(\serial_flash_inf_cmd_gen_inst|Selector9~4_combout ),
	.Selector17(\serial_flash_inf_cmd_gen_inst|Selector17~0_combout ),
	.mem_addr_reg_6(\xip_controller|mem_addr_reg[6]~q ),
	.mem_addr_reg_14(\xip_controller|mem_addr_reg[14]~q ),
	.addr_bytes_xip_0(\xip_controller|addr_bytes_xip[0]~0_combout ),
	.mem_addr_reg_10(\xip_controller|mem_addr_reg[10]~q ),
	.mem_addr_reg_18(\xip_controller|mem_addr_reg[18]~q ),
	.mem_addr_reg_2(\xip_controller|mem_addr_reg[2]~q ),
	.mem_addr_reg_8(\xip_controller|mem_addr_reg[8]~q ),
	.mem_addr_reg_16(\xip_controller|mem_addr_reg[16]~q ),
	.mem_addr_reg_0(\xip_controller|mem_addr_reg[0]~q ),
	.mem_addr_reg_15(\xip_controller|mem_addr_reg[15]~q ),
	.mem_addr_reg_7(\xip_controller|mem_addr_reg[7]~q ),
	.WideOr19(\xip_controller|WideOr19~0_combout ),
	.mem_addr_reg_17(\xip_controller|mem_addr_reg[17]~q ),
	.mem_addr_reg_9(\xip_controller|mem_addr_reg[9]~q ),
	.mem_addr_reg_1(\xip_controller|mem_addr_reg[1]~q ),
	.mem_addr_reg_19(\xip_controller|mem_addr_reg[19]~q ),
	.mem_addr_reg_11(\xip_controller|mem_addr_reg[11]~q ),
	.mem_addr_reg_3(\xip_controller|mem_addr_reg[3]~q ),
	.mem_addr_reg_12(\xip_controller|mem_addr_reg[12]~q ),
	.mem_addr_reg_20(\xip_controller|mem_addr_reg[20]~q ),
	.mem_addr_reg_4(\xip_controller|mem_addr_reg[4]~q ),
	.mem_addr_reg_13(\xip_controller|mem_addr_reg[13]~q ),
	.mem_addr_reg_5(\xip_controller|mem_addr_reg[5]~q ),
	.has_dummy(\csr_controller|has_dummy~q ),
	.cmd_data_12(\xip_controller|cmd_data[12]~combout ),
	.out_payload_31(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[31]~q ),
	.clk_clk(clk_clk));

flashLoader_flashLoader_intel_generic_serial_flash_interface_top_0_multiplexer multiplexer(
	.stateST_IDLE(\csr_controller|state.ST_IDLE~q ),
	.csr_flash_cmd_wr_data_0_data_0(\csr_controller|csr_flash_cmd_wr_data_0_data[0]~q ),
	.csr_flash_cmd_wr_data_1_data_0(\csr_controller|csr_flash_cmd_wr_data_1_data[0]~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.csr_flash_cmd_wr_data_0_data_1(\csr_controller|csr_flash_cmd_wr_data_0_data[1]~q ),
	.csr_flash_cmd_wr_data_1_data_1(\csr_controller|csr_flash_cmd_wr_data_1_data[1]~q ),
	.csr_flash_cmd_wr_data_0_data_2(\csr_controller|csr_flash_cmd_wr_data_0_data[2]~q ),
	.csr_flash_cmd_wr_data_1_data_2(\csr_controller|csr_flash_cmd_wr_data_1_data[2]~q ),
	.csr_flash_cmd_wr_data_0_data_3(\csr_controller|csr_flash_cmd_wr_data_0_data[3]~q ),
	.csr_flash_cmd_wr_data_1_data_3(\csr_controller|csr_flash_cmd_wr_data_1_data[3]~q ),
	.csr_control_data_4(\csr_controller|csr_control_data[4]~q ),
	.csr_flash_cmd_wr_data_1_data_4(\csr_controller|csr_flash_cmd_wr_data_1_data[4]~q ),
	.csr_flash_cmd_wr_data_0_data_4(\csr_controller|csr_flash_cmd_wr_data_0_data[4]~q ),
	.csr_control_data_5(\csr_controller|csr_control_data[5]~q ),
	.csr_flash_cmd_wr_data_1_data_5(\csr_controller|csr_flash_cmd_wr_data_1_data[5]~q ),
	.csr_flash_cmd_wr_data_0_data_5(\csr_controller|csr_flash_cmd_wr_data_0_data[5]~q ),
	.csr_control_data_6(\csr_controller|csr_control_data[6]~q ),
	.csr_flash_cmd_wr_data_1_data_6(\csr_controller|csr_flash_cmd_wr_data_1_data[6]~q ),
	.csr_flash_cmd_wr_data_0_data_6(\csr_controller|csr_flash_cmd_wr_data_0_data[6]~q ),
	.csr_control_data_7(\csr_controller|csr_control_data[7]~q ),
	.csr_flash_cmd_wr_data_1_data_7(\csr_controller|csr_flash_cmd_wr_data_1_data[7]~q ),
	.csr_flash_cmd_wr_data_0_data_7(\csr_controller|csr_flash_cmd_wr_data_0_data[7]~q ),
	.csr_flash_cmd_wr_data_0_data_8(\csr_controller|csr_flash_cmd_wr_data_0_data[8]~q ),
	.csr_flash_cmd_wr_data_1_data_8(\csr_controller|csr_flash_cmd_wr_data_1_data[8]~q ),
	.csr_flash_cmd_wr_data_0_data_9(\csr_controller|csr_flash_cmd_wr_data_0_data[9]~q ),
	.csr_flash_cmd_wr_data_1_data_9(\csr_controller|csr_flash_cmd_wr_data_1_data[9]~q ),
	.csr_flash_cmd_wr_data_0_data_10(\csr_controller|csr_flash_cmd_wr_data_0_data[10]~q ),
	.csr_flash_cmd_wr_data_1_data_10(\csr_controller|csr_flash_cmd_wr_data_1_data[10]~q ),
	.csr_rd_inst_data_11(\csr_controller|csr_rd_inst_data[11]~q ),
	.csr_flash_cmd_wr_data_0_data_11(\csr_controller|csr_flash_cmd_wr_data_0_data[11]~q ),
	.csr_flash_cmd_wr_data_1_data_11(\csr_controller|csr_flash_cmd_wr_data_1_data[11]~q ),
	.csr_rd_inst_data_12(\csr_controller|csr_rd_inst_data[12]~q ),
	.csr_flash_cmd_wr_data_0_data_13(\csr_controller|csr_flash_cmd_wr_data_0_data[13]~q ),
	.csr_flash_cmd_wr_data_1_data_13(\csr_controller|csr_flash_cmd_wr_data_1_data[13]~q ),
	.csr_flash_cmd_wr_data_0_data_14(\csr_controller|csr_flash_cmd_wr_data_0_data[14]~q ),
	.csr_flash_cmd_wr_data_1_data_14(\csr_controller|csr_flash_cmd_wr_data_1_data[14]~q ),
	.csr_flash_cmd_wr_data_0_data_15(\csr_controller|csr_flash_cmd_wr_data_0_data[15]~q ),
	.csr_flash_cmd_wr_data_1_data_15(\csr_controller|csr_flash_cmd_wr_data_1_data[15]~q ),
	.csr_flash_cmd_wr_data_0_data_16(\csr_controller|csr_flash_cmd_wr_data_0_data[16]~q ),
	.csr_flash_cmd_wr_data_1_data_16(\csr_controller|csr_flash_cmd_wr_data_1_data[16]~q ),
	.csr_flash_cmd_wr_data_0_data_17(\csr_controller|csr_flash_cmd_wr_data_0_data[17]~q ),
	.csr_flash_cmd_wr_data_1_data_17(\csr_controller|csr_flash_cmd_wr_data_1_data[17]~q ),
	.csr_flash_cmd_wr_data_0_data_18(\csr_controller|csr_flash_cmd_wr_data_0_data[18]~q ),
	.csr_flash_cmd_wr_data_1_data_18(\csr_controller|csr_flash_cmd_wr_data_1_data[18]~q ),
	.csr_flash_cmd_wr_data_0_data_19(\csr_controller|csr_flash_cmd_wr_data_0_data[19]~q ),
	.csr_flash_cmd_wr_data_1_data_19(\csr_controller|csr_flash_cmd_wr_data_1_data[19]~q ),
	.csr_flash_cmd_wr_data_0_data_20(\csr_controller|csr_flash_cmd_wr_data_0_data[20]~q ),
	.csr_flash_cmd_wr_data_1_data_20(\csr_controller|csr_flash_cmd_wr_data_1_data[20]~q ),
	.csr_flash_cmd_wr_data_0_data_21(\csr_controller|csr_flash_cmd_wr_data_0_data[21]~q ),
	.csr_flash_cmd_wr_data_1_data_21(\csr_controller|csr_flash_cmd_wr_data_1_data[21]~q ),
	.csr_flash_cmd_wr_data_0_data_22(\csr_controller|csr_flash_cmd_wr_data_0_data[22]~q ),
	.csr_flash_cmd_wr_data_1_data_22(\csr_controller|csr_flash_cmd_wr_data_1_data[22]~q ),
	.csr_flash_cmd_wr_data_0_data_23(\csr_controller|csr_flash_cmd_wr_data_0_data[23]~q ),
	.csr_flash_cmd_wr_data_1_data_23(\csr_controller|csr_flash_cmd_wr_data_1_data[23]~q ),
	.csr_flash_cmd_wr_data_0_data_24(\csr_controller|csr_flash_cmd_wr_data_0_data[24]~q ),
	.csr_flash_cmd_wr_data_1_data_24(\csr_controller|csr_flash_cmd_wr_data_1_data[24]~q ),
	.csr_flash_cmd_wr_data_0_data_25(\csr_controller|csr_flash_cmd_wr_data_0_data[25]~q ),
	.csr_flash_cmd_wr_data_1_data_25(\csr_controller|csr_flash_cmd_wr_data_1_data[25]~q ),
	.csr_flash_cmd_wr_data_0_data_26(\csr_controller|csr_flash_cmd_wr_data_0_data[26]~q ),
	.csr_flash_cmd_wr_data_1_data_26(\csr_controller|csr_flash_cmd_wr_data_1_data[26]~q ),
	.csr_flash_cmd_wr_data_0_data_27(\csr_controller|csr_flash_cmd_wr_data_0_data[27]~q ),
	.csr_flash_cmd_wr_data_1_data_27(\csr_controller|csr_flash_cmd_wr_data_1_data[27]~q ),
	.csr_flash_cmd_wr_data_0_data_28(\csr_controller|csr_flash_cmd_wr_data_0_data[28]~q ),
	.csr_flash_cmd_wr_data_1_data_28(\csr_controller|csr_flash_cmd_wr_data_1_data[28]~q ),
	.csr_flash_cmd_wr_data_0_data_29(\csr_controller|csr_flash_cmd_wr_data_0_data[29]~q ),
	.csr_flash_cmd_wr_data_1_data_29(\csr_controller|csr_flash_cmd_wr_data_1_data[29]~q ),
	.csr_flash_cmd_wr_data_0_data_30(\csr_controller|csr_flash_cmd_wr_data_0_data[30]~q ),
	.csr_flash_cmd_wr_data_1_data_30(\csr_controller|csr_flash_cmd_wr_data_1_data[30]~q ),
	.stateST_WAIT_RSP(\csr_controller|state.ST_WAIT_RSP~q ),
	.saved_grant_1(\multiplexer|saved_grant[1]~q ),
	.stateST_SEND_HEADER(\csr_controller|state.ST_SEND_HEADER~q ),
	.saved_grant_0(\multiplexer|saved_grant[0]~q ),
	.current_stateSTATE_WR_CMD(\xip_controller|current_state.STATE_WR_CMD~q ),
	.current_stateSTATE_STATUS_CMD(\xip_controller|current_state.STATE_STATUS_CMD~q ),
	.current_stateSTATE_POLL_CMD(\xip_controller|current_state.STATE_POLL_CMD~q ),
	.current_stateSTATE_READ_CMD(\xip_controller|current_state.STATE_READ_CMD~q ),
	.WideOr13(\xip_controller|WideOr13~0_combout ),
	.src_startofpacket1(\multiplexer|src_startofpacket~combout ),
	.src_valid(\multiplexer|src_valid~0_combout ),
	.current_stateSTATE_WR_DATA(\xip_controller|current_state.STATE_WR_DATA~q ),
	.cmd_valid(\xip_controller|cmd_valid~0_combout ),
	.stateST_SEND_DATA(\serial_flash_inf_cmd_gen_inst|state.ST_SEND_DATA~q ),
	.Selector18(\serial_flash_inf_cmd_gen_inst|Selector18~2_combout ),
	.WideOr0(\qspi_inf_inst|demultiplexer_inst|WideOr0~3_combout ),
	.in_ready(\qspi_inf_inst|adapter_8_4_inst|in_ready~combout ),
	.WideOr01(\qspi_inf_inst|demultiplexer_inst|WideOr0~4_combout ),
	.adap_out_cmd_ready(\serial_flash_inf_cmd_gen_inst|adap_out_cmd_ready~0_combout ),
	.Selector181(\serial_flash_inf_cmd_gen_inst|Selector18~3_combout ),
	.stateST_SEND_DATA_1(\csr_controller|state.ST_SEND_DATA_1~q ),
	.stateST_SEND_DATA_0(\csr_controller|state.ST_SEND_DATA_0~q ),
	.has_data_in(\csr_controller|has_data_in~q ),
	.more_than_4bytes_data(\csr_controller|more_than_4bytes_data~q ),
	.src_payload_0(\multiplexer|src_payload[0]~1_combout ),
	.Selector182(\serial_flash_inf_cmd_gen_inst|Selector18~5_combout ),
	.sink0_ready(\multiplexer|sink0_ready~1_combout ),
	.src_data_30(\multiplexer|src_data[30]~3_combout ),
	.is_burst_reg(\xip_controller|is_burst_reg~q ),
	.mem_write_data_reg_30(\xip_controller|mem_write_data_reg[30]~q ),
	.mem_byteenable_reg_0(\xip_controller|mem_byteenable_reg[0]~q ),
	.mem_byteenable_reg_3(\xip_controller|mem_byteenable_reg[3]~q ),
	.mem_byteenable_reg_2(\xip_controller|mem_byteenable_reg[2]~q ),
	.mem_byteenable_reg_1(\xip_controller|mem_byteenable_reg[1]~q ),
	.src_data_301(\multiplexer|src_data[30]~5_combout ),
	.out_payload_30(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[30]~q ),
	.cmd_valid1(\xip_controller|cmd_valid~1_combout ),
	.src_data_302(\multiplexer|src_data[30]~7_combout ),
	.src_data_303(\multiplexer|src_data[30]~8_combout ),
	.src_data_29(\multiplexer|src_data[29]~10_combout ),
	.mem_write_data_reg_29(\xip_controller|mem_write_data_reg[29]~q ),
	.out_payload_29(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[29]~q ),
	.src_data_291(\multiplexer|src_data[29]~12_combout ),
	.src_data_292(\multiplexer|src_data[29]~13_combout ),
	.src_data_28(\multiplexer|src_data[28]~15_combout ),
	.mem_write_data_reg_28(\xip_controller|mem_write_data_reg[28]~q ),
	.out_payload_28(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[28]~q ),
	.src_data_281(\multiplexer|src_data[28]~17_combout ),
	.src_data_282(\multiplexer|src_data[28]~18_combout ),
	.src_data_27(\multiplexer|src_data[27]~20_combout ),
	.mem_write_data_reg_27(\xip_controller|mem_write_data_reg[27]~q ),
	.out_payload_27(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[27]~q ),
	.src_data_271(\multiplexer|src_data[27]~22_combout ),
	.src_data_272(\multiplexer|src_data[27]~23_combout ),
	.WideOr11(\multiplexer|WideOr1~combout ),
	.out_payload_32(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[32]~q ),
	.src_payload_01(\multiplexer|src_payload[0]~3_combout ),
	.sink1_ready1(\multiplexer|sink1_ready~combout ),
	.Selector34(\csr_controller|Selector34~0_combout ),
	.has_data_out(\csr_controller|has_data_out~q ),
	.src_data_11(\multiplexer|src_data[11]~25_combout ),
	.cmd_data_11(\xip_controller|cmd_data[11]~combout ),
	.src_data_111(\multiplexer|src_data[11]~26_combout ),
	.numb_data_0(\csr_controller|numb_data[0]~q ),
	.Add1(\xip_controller|Add1~1_combout ),
	.Selector20(\xip_controller|Selector20~0_combout ),
	.out_payload_18(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[18]~q ),
	.mem_write_data_reg_18(\xip_controller|mem_write_data_reg[18]~q ),
	.src_data_18(\multiplexer|src_data[18]~32_combout ),
	.numb_data_1(\csr_controller|numb_data[1]~q ),
	.src_data_19(\multiplexer|src_data[19]~34_combout ),
	.Add11(\xip_controller|Add1~2_combout ),
	.mem_write_data_reg_19(\xip_controller|mem_write_data_reg[19]~q ),
	.out_payload_19(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[19]~q ),
	.src_data_191(\multiplexer|src_data[19]~37_combout ),
	.src_data_192(\multiplexer|src_data[19]~38_combout ),
	.numb_data_3(\csr_controller|numb_data[3]~q ),
	.src_data_21(\multiplexer|src_data[21]~40_combout ),
	.mem_write_data_reg_21(\xip_controller|mem_write_data_reg[21]~q ),
	.out_payload_21(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[21]~q ),
	.mem_burstcount_reg_1(\xip_controller|mem_burstcount_reg[1]~q ),
	.src_data_211(\multiplexer|src_data[21]~43_combout ),
	.src_data_212(\multiplexer|src_data[21]~44_combout ),
	.numb_data_2(\csr_controller|numb_data[2]~q ),
	.src_data_20(\multiplexer|src_data[20]~46_combout ),
	.mem_write_data_reg_20(\xip_controller|mem_write_data_reg[20]~q ),
	.out_payload_20(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[20]~q ),
	.mem_burstcount_reg_0(\xip_controller|mem_burstcount_reg[0]~q ),
	.src_data_201(\multiplexer|src_data[20]~50_combout ),
	.src_data_202(\multiplexer|src_data[20]~51_combout ),
	.mem_write_data_reg_22(\xip_controller|mem_write_data_reg[22]~q ),
	.out_payload_22(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[22]~q ),
	.mem_burstcount_reg_2(\xip_controller|mem_burstcount_reg[2]~q ),
	.src_data_22(\multiplexer|src_data[22]~55_combout ),
	.mem_write_data_reg_23(\xip_controller|mem_write_data_reg[23]~q ),
	.out_payload_23(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[23]~q ),
	.mem_burstcount_reg_3(\xip_controller|mem_burstcount_reg[3]~q ),
	.src_data_23(\multiplexer|src_data[23]~59_combout ),
	.mem_write_data_reg_24(\xip_controller|mem_write_data_reg[24]~q ),
	.out_payload_24(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[24]~q ),
	.mem_burstcount_reg_4(\xip_controller|mem_burstcount_reg[4]~q ),
	.src_data_24(\multiplexer|src_data[24]~63_combout ),
	.mem_write_data_reg_25(\xip_controller|mem_write_data_reg[25]~q ),
	.out_payload_25(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[25]~q ),
	.mem_burstcount_reg_5(\xip_controller|mem_burstcount_reg[5]~q ),
	.src_data_25(\multiplexer|src_data[25]~67_combout ),
	.mem_write_data_reg_26(\xip_controller|mem_write_data_reg[26]~q ),
	.out_payload_26(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[26]~q ),
	.mem_burstcount_reg_6(\xip_controller|mem_burstcount_reg[6]~q ),
	.src_data_26(\multiplexer|src_data[26]~71_combout ),
	.src_data_10(\multiplexer|src_data[10]~73_combout ),
	.cmd_data_10(\xip_controller|cmd_data[10]~combout ),
	.src_data_101(\multiplexer|src_data[10]~74_combout ),
	.has_addr(\csr_controller|has_addr~q ),
	.src_data_8(\multiplexer|src_data[8]~76_combout ),
	.cmd_data_8(\xip_controller|cmd_data[8]~combout ),
	.src_data_81(\multiplexer|src_data[8]~77_combout ),
	.numb_dummy_0(\csr_controller|numb_dummy[0]~q ),
	.src_data_13(\multiplexer|src_data[13]~79_combout ),
	.cmd_data_13(\xip_controller|cmd_data[13]~combout ),
	.src_data_131(\multiplexer|src_data[13]~80_combout ),
	.numb_dummy_4(\csr_controller|numb_dummy[4]~q ),
	.src_data_17(\multiplexer|src_data[17]~82_combout ),
	.mem_write_data_reg_17(\xip_controller|mem_write_data_reg[17]~q ),
	.out_payload_17(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[17]~q ),
	.src_data_171(\multiplexer|src_data[17]~84_combout ),
	.src_data_172(\multiplexer|src_data[17]~85_combout ),
	.numb_dummy_3(\csr_controller|numb_dummy[3]~q ),
	.src_data_16(\multiplexer|src_data[16]~87_combout ),
	.mem_write_data_reg_16(\xip_controller|mem_write_data_reg[16]~q ),
	.out_payload_16(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[16]~q ),
	.src_data_161(\multiplexer|src_data[16]~89_combout ),
	.src_data_162(\multiplexer|src_data[16]~90_combout ),
	.numb_dummy_2(\csr_controller|numb_dummy[2]~q ),
	.src_data_15(\multiplexer|src_data[15]~92_combout ),
	.cmd_data_15(\xip_controller|cmd_data[15]~combout ),
	.src_data_151(\multiplexer|src_data[15]~93_combout ),
	.numb_dummy_1(\csr_controller|numb_dummy[1]~q ),
	.src_data_14(\multiplexer|src_data[14]~95_combout ),
	.cmd_data_14(\xip_controller|cmd_data[14]~combout ),
	.src_data_141(\multiplexer|src_data[14]~96_combout ),
	.is_4bytes_addr(\csr_controller|is_4bytes_addr~q ),
	.src_data_9(\multiplexer|src_data[9]~98_combout ),
	.cmd_data_9(\xip_controller|cmd_data[9]~combout ),
	.src_data_91(\multiplexer|src_data[9]~99_combout ),
	.opcode_0(\csr_controller|opcode[0]~q ),
	.out_payload_0(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[0]~q ),
	.cmd_data_0(\xip_controller|cmd_data[0]~36_combout ),
	.src_data_0(\multiplexer|src_data[0]~102_combout ),
	.opcode_4(\csr_controller|opcode[4]~q ),
	.out_payload_4(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[4]~q ),
	.cmd_data_4(\xip_controller|cmd_data[4]~43_combout ),
	.src_data_4(\multiplexer|src_data[4]~105_combout ),
	.opcode_2(\csr_controller|opcode[2]~q ),
	.out_payload_2(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[2]~q ),
	.cmd_data_2(\xip_controller|cmd_data[2]~50_combout ),
	.src_data_2(\multiplexer|src_data[2]~108_combout ),
	.opcode_1(\csr_controller|opcode[1]~q ),
	.out_payload_1(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[1]~q ),
	.cmd_data_1(\xip_controller|cmd_data[1]~57_combout ),
	.src_data_1(\multiplexer|src_data[1]~111_combout ),
	.opcode_3(\csr_controller|opcode[3]~q ),
	.out_payload_3(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[3]~q ),
	.cmd_data_3(\xip_controller|cmd_data[3]~64_combout ),
	.src_data_3(\multiplexer|src_data[3]~114_combout ),
	.opcode_5(\csr_controller|opcode[5]~q ),
	.out_payload_5(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[5]~q ),
	.cmd_data_5(\xip_controller|cmd_data[5]~71_combout ),
	.src_data_5(\multiplexer|src_data[5]~117_combout ),
	.opcode_6(\csr_controller|opcode[6]~q ),
	.out_payload_6(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[6]~q ),
	.cmd_data_6(\xip_controller|cmd_data[6]~78_combout ),
	.src_data_6(\multiplexer|src_data[6]~120_combout ),
	.opcode_7(\csr_controller|opcode[7]~q ),
	.out_payload_7(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[7]~q ),
	.cmd_data_7(\xip_controller|cmd_data[7]~85_combout ),
	.src_data_7(\multiplexer|src_data[7]~123_combout ),
	.clk_clk(clk_clk));

flashLoader_flashLoader_intel_generic_serial_flash_interface_top_0_merlin_demultiplexer_0 merlin_demultiplexer_0(
	.in_cmd_channel_reg_1(\serial_flash_inf_cmd_gen_inst|in_cmd_channel_reg[1]~q ),
	.stateST_WAIT_RSP(\csr_controller|state.ST_WAIT_RSP~q ),
	.sink_ready(\merlin_demultiplexer_0|sink_ready~0_combout ),
	.in_cmd_channel_reg_0(\serial_flash_inf_cmd_gen_inst|in_cmd_channel_reg[0]~q ),
	.WideOr01(\merlin_demultiplexer_0|WideOr0~combout ));

flashLoader_flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller xip_controller(
	.hold_waitrequest1(\xip_controller|hold_waitrequest~q ),
	.mem_waitrequest(mem_waitrequest),
	.mem_rddata_0(mem_rddata_0),
	.mem_rddata_1(mem_rddata_1),
	.mem_rddata_2(mem_rddata_2),
	.mem_rddata_3(mem_rddata_3),
	.mem_rddata_4(mem_rddata_4),
	.mem_rddata_5(mem_rddata_5),
	.mem_rddata_6(mem_rddata_6),
	.mem_rddata_7(mem_rddata_7),
	.mem_rddata_8(mem_rddata_8),
	.mem_rddata_9(mem_rddata_9),
	.mem_rddata_10(mem_rddata_10),
	.mem_rddata_11(mem_rddata_11),
	.mem_rddata_12(mem_rddata_12),
	.mem_rddata_13(mem_rddata_13),
	.mem_rddata_14(mem_rddata_14),
	.mem_rddata_15(mem_rddata_15),
	.mem_rddata_16(mem_rddata_16),
	.mem_rddata_17(mem_rddata_17),
	.mem_rddata_18(mem_rddata_18),
	.mem_rddata_19(mem_rddata_19),
	.mem_rddata_20(mem_rddata_20),
	.mem_rddata_21(mem_rddata_21),
	.mem_rddata_22(mem_rddata_22),
	.mem_rddata_23(mem_rddata_23),
	.mem_rddata_24(mem_rddata_24),
	.mem_rddata_25(mem_rddata_25),
	.mem_rddata_26(mem_rddata_26),
	.mem_rddata_27(mem_rddata_27),
	.mem_rddata_28(mem_rddata_28),
	.mem_rddata_29(mem_rddata_29),
	.mem_rddata_30(mem_rddata_30),
	.mem_rddata_31(mem_rddata_31),
	.mem_rddatavalid1(mem_rddatavalid),
	.csr_wr_inst_data_0(\csr_controller|csr_wr_inst_data[0]~q ),
	.csr_rd_inst_data_0(\csr_controller|csr_rd_inst_data[0]~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.csr_wr_inst_data_1(\csr_controller|csr_wr_inst_data[1]~q ),
	.csr_rd_inst_data_1(\csr_controller|csr_rd_inst_data[1]~q ),
	.csr_wr_inst_data_2(\csr_controller|csr_wr_inst_data[2]~q ),
	.csr_rd_inst_data_2(\csr_controller|csr_rd_inst_data[2]~q ),
	.csr_wr_inst_data_3(\csr_controller|csr_wr_inst_data[3]~q ),
	.csr_rd_inst_data_3(\csr_controller|csr_rd_inst_data[3]~q ),
	.csr_wr_inst_data_4(\csr_controller|csr_wr_inst_data[4]~q ),
	.csr_rd_inst_data_4(\csr_controller|csr_rd_inst_data[4]~q ),
	.csr_wr_inst_data_5(\csr_controller|csr_wr_inst_data[5]~q ),
	.csr_rd_inst_data_5(\csr_controller|csr_rd_inst_data[5]~q ),
	.csr_wr_inst_data_6(\csr_controller|csr_wr_inst_data[6]~q ),
	.csr_rd_inst_data_6(\csr_controller|csr_rd_inst_data[6]~q ),
	.csr_wr_inst_data_7(\csr_controller|csr_wr_inst_data[7]~q ),
	.csr_rd_inst_data_7(\csr_controller|csr_rd_inst_data[7]~q ),
	.csr_rd_inst_data_8(\csr_controller|csr_rd_inst_data[8]~q ),
	.csr_control_data_8(\csr_controller|csr_control_data[8]~q ),
	.csr_wr_inst_data_8(\csr_controller|csr_wr_inst_data[8]~q ),
	.csr_rd_inst_data_9(\csr_controller|csr_rd_inst_data[9]~q ),
	.csr_wr_inst_data_9(\csr_controller|csr_wr_inst_data[9]~q ),
	.csr_rd_inst_data_10(\csr_controller|csr_rd_inst_data[10]~q ),
	.csr_wr_inst_data_10(\csr_controller|csr_wr_inst_data[10]~q ),
	.csr_rd_inst_data_11(\csr_controller|csr_rd_inst_data[11]~q ),
	.csr_wr_inst_data_11(\csr_controller|csr_wr_inst_data[11]~q ),
	.csr_rd_inst_data_12(\csr_controller|csr_rd_inst_data[12]~q ),
	.csr_wr_inst_data_12(\csr_controller|csr_wr_inst_data[12]~q ),
	.csr_wr_inst_data_13(\csr_controller|csr_wr_inst_data[13]~q ),
	.csr_wr_inst_data_14(\csr_controller|csr_wr_inst_data[14]~q ),
	.csr_wr_inst_data_15(\csr_controller|csr_wr_inst_data[15]~q ),
	.stateST_SEND_DUMMY_RSP(\serial_flash_inf_cmd_gen_inst|state.ST_SEND_DUMMY_RSP~q ),
	.out_valid(\serial_flash_inf_cmd_gen_inst|data_adapter_8_32_inst|out_valid~q ),
	.out_endofpacket(\serial_flash_inf_cmd_gen_inst|data_adapter_8_32_inst|out_endofpacket~q ),
	.out_data_0(\serial_flash_inf_cmd_gen_inst|data_adapter_8_32_inst|out_data[0]~q ),
	.out_rsp_data_0(\serial_flash_inf_cmd_gen_inst|out_rsp_data[0]~0_combout ),
	.current_stateSTATE_READ_DATA(\xip_controller|current_state.STATE_READ_DATA~q ),
	.out_rsp_data_1(\serial_flash_inf_cmd_gen_inst|out_rsp_data[1]~1_combout ),
	.out_rsp_data_2(\serial_flash_inf_cmd_gen_inst|out_rsp_data[2]~2_combout ),
	.out_rsp_data_3(\serial_flash_inf_cmd_gen_inst|out_rsp_data[3]~3_combout ),
	.out_rsp_data_4(\serial_flash_inf_cmd_gen_inst|out_rsp_data[4]~4_combout ),
	.out_rsp_data_5(\serial_flash_inf_cmd_gen_inst|out_rsp_data[5]~5_combout ),
	.out_rsp_data_6(\serial_flash_inf_cmd_gen_inst|out_rsp_data[6]~6_combout ),
	.out_rsp_data_7(\serial_flash_inf_cmd_gen_inst|out_rsp_data[7]~7_combout ),
	.out_rsp_data_8(\serial_flash_inf_cmd_gen_inst|out_rsp_data[8]~8_combout ),
	.out_rsp_data_9(\serial_flash_inf_cmd_gen_inst|out_rsp_data[9]~9_combout ),
	.out_rsp_data_10(\serial_flash_inf_cmd_gen_inst|out_rsp_data[10]~10_combout ),
	.out_rsp_data_11(\serial_flash_inf_cmd_gen_inst|out_rsp_data[11]~11_combout ),
	.out_rsp_data_12(\serial_flash_inf_cmd_gen_inst|out_rsp_data[12]~12_combout ),
	.out_rsp_data_13(\serial_flash_inf_cmd_gen_inst|out_rsp_data[13]~13_combout ),
	.out_rsp_data_14(\serial_flash_inf_cmd_gen_inst|out_rsp_data[14]~14_combout ),
	.out_rsp_data_15(\serial_flash_inf_cmd_gen_inst|out_rsp_data[15]~15_combout ),
	.out_rsp_data_16(\serial_flash_inf_cmd_gen_inst|out_rsp_data[16]~16_combout ),
	.out_rsp_data_17(\serial_flash_inf_cmd_gen_inst|out_rsp_data[17]~17_combout ),
	.out_rsp_data_18(\serial_flash_inf_cmd_gen_inst|out_rsp_data[18]~18_combout ),
	.out_rsp_data_19(\serial_flash_inf_cmd_gen_inst|out_rsp_data[19]~19_combout ),
	.out_rsp_data_20(\serial_flash_inf_cmd_gen_inst|out_rsp_data[20]~20_combout ),
	.out_rsp_data_21(\serial_flash_inf_cmd_gen_inst|out_rsp_data[21]~21_combout ),
	.out_rsp_data_22(\serial_flash_inf_cmd_gen_inst|out_rsp_data[22]~22_combout ),
	.out_rsp_data_23(\serial_flash_inf_cmd_gen_inst|out_rsp_data[23]~23_combout ),
	.out_rsp_data_24(\serial_flash_inf_cmd_gen_inst|out_rsp_data[24]~24_combout ),
	.out_rsp_data_25(\serial_flash_inf_cmd_gen_inst|out_rsp_data[25]~25_combout ),
	.out_rsp_data_26(\serial_flash_inf_cmd_gen_inst|out_rsp_data[26]~26_combout ),
	.out_rsp_data_27(\serial_flash_inf_cmd_gen_inst|out_rsp_data[27]~27_combout ),
	.out_rsp_data_28(\serial_flash_inf_cmd_gen_inst|out_rsp_data[28]~28_combout ),
	.out_rsp_data_29(\serial_flash_inf_cmd_gen_inst|out_rsp_data[29]~29_combout ),
	.out_rsp_data_30(\serial_flash_inf_cmd_gen_inst|out_rsp_data[30]~30_combout ),
	.out_rsp_data_31(\serial_flash_inf_cmd_gen_inst|out_rsp_data[31]~31_combout ),
	.in_cmd_channel_reg_0(\serial_flash_inf_cmd_gen_inst|in_cmd_channel_reg[0]~q ),
	.saved_grant_0(\multiplexer|saved_grant[0]~q ),
	.current_stateSTATE_WR_CMD(\xip_controller|current_state.STATE_WR_CMD~q ),
	.current_stateSTATE_STATUS_CMD(\xip_controller|current_state.STATE_STATUS_CMD~q ),
	.current_stateSTATE_POLL_CMD(\xip_controller|current_state.STATE_POLL_CMD~q ),
	.current_stateSTATE_READ_CMD(\xip_controller|current_state.STATE_READ_CMD~q ),
	.WideOr13(\xip_controller|WideOr13~0_combout ),
	.current_stateSTATE_WR_DATA(\xip_controller|current_state.STATE_WR_DATA~q ),
	.cmd_valid(\xip_controller|cmd_valid~0_combout ),
	.Selector18(\serial_flash_inf_cmd_gen_inst|Selector18~2_combout ),
	.adap_out_cmd_ready(\serial_flash_inf_cmd_gen_inst|adap_out_cmd_ready~0_combout ),
	.Selector181(\serial_flash_inf_cmd_gen_inst|Selector18~3_combout ),
	.sink0_ready(\multiplexer|sink0_ready~1_combout ),
	.is_burst_reg1(\xip_controller|is_burst_reg~q ),
	.mem_write_data_reg_30(\xip_controller|mem_write_data_reg[30]~q ),
	.mem_byteenable_reg_0(\xip_controller|mem_byteenable_reg[0]~q ),
	.mem_byteenable_reg_3(\xip_controller|mem_byteenable_reg[3]~q ),
	.mem_byteenable_reg_2(\xip_controller|mem_byteenable_reg[2]~q ),
	.mem_byteenable_reg_1(\xip_controller|mem_byteenable_reg[1]~q ),
	.out_payload_30(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[30]~q ),
	.cmd_valid1(\xip_controller|cmd_valid~1_combout ),
	.mem_write_data_reg_29(\xip_controller|mem_write_data_reg[29]~q ),
	.out_payload_29(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[29]~q ),
	.mem_write_data_reg_28(\xip_controller|mem_write_data_reg[28]~q ),
	.out_payload_28(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[28]~q ),
	.mem_write_data_reg_27(\xip_controller|mem_write_data_reg[27]~q ),
	.out_payload_27(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[27]~q ),
	.out_payload_32(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[32]~q ),
	.cmd_data_11(\xip_controller|cmd_data[11]~combout ),
	.Add1(\xip_controller|Add1~1_combout ),
	.Selector20(\xip_controller|Selector20~0_combout ),
	.out_payload_18(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[18]~q ),
	.mem_write_data_reg_18(\xip_controller|mem_write_data_reg[18]~q ),
	.Add11(\xip_controller|Add1~2_combout ),
	.mem_write_data_reg_19(\xip_controller|mem_write_data_reg[19]~q ),
	.out_payload_19(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[19]~q ),
	.mem_write_data_reg_21(\xip_controller|mem_write_data_reg[21]~q ),
	.out_payload_21(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[21]~q ),
	.mem_burstcount_reg_1(\xip_controller|mem_burstcount_reg[1]~q ),
	.mem_write_data_reg_20(\xip_controller|mem_write_data_reg[20]~q ),
	.out_payload_20(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[20]~q ),
	.mem_burstcount_reg_0(\xip_controller|mem_burstcount_reg[0]~q ),
	.mem_write_data_reg_22(\xip_controller|mem_write_data_reg[22]~q ),
	.out_payload_22(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[22]~q ),
	.mem_burstcount_reg_2(\xip_controller|mem_burstcount_reg[2]~q ),
	.mem_write_data_reg_23(\xip_controller|mem_write_data_reg[23]~q ),
	.out_payload_23(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[23]~q ),
	.mem_burstcount_reg_3(\xip_controller|mem_burstcount_reg[3]~q ),
	.mem_write_data_reg_24(\xip_controller|mem_write_data_reg[24]~q ),
	.out_payload_24(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[24]~q ),
	.mem_burstcount_reg_4(\xip_controller|mem_burstcount_reg[4]~q ),
	.mem_write_data_reg_25(\xip_controller|mem_write_data_reg[25]~q ),
	.out_payload_25(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[25]~q ),
	.mem_burstcount_reg_5(\xip_controller|mem_burstcount_reg[5]~q ),
	.mem_write_data_reg_26(\xip_controller|mem_write_data_reg[26]~q ),
	.out_payload_26(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[26]~q ),
	.mem_burstcount_reg_6(\xip_controller|mem_burstcount_reg[6]~q ),
	.cmd_data_10(\xip_controller|cmd_data[10]~combout ),
	.cmd_data_8(\xip_controller|cmd_data[8]~combout ),
	.cmd_data_13(\xip_controller|cmd_data[13]~combout ),
	.mem_write_data_reg_17(\xip_controller|mem_write_data_reg[17]~q ),
	.out_payload_17(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[17]~q ),
	.mem_write_data_reg_16(\xip_controller|mem_write_data_reg[16]~q ),
	.out_payload_16(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[16]~q ),
	.mem_write_data_reg_31(\xip_controller|mem_write_data_reg[31]~q ),
	.cmd_data_15(\xip_controller|cmd_data[15]~combout ),
	.cmd_data_14(\xip_controller|cmd_data[14]~combout ),
	.cmd_data_9(\xip_controller|cmd_data[9]~combout ),
	.mem_addr_reg_6(\xip_controller|mem_addr_reg[6]~q ),
	.mem_addr_reg_14(\xip_controller|mem_addr_reg[14]~q ),
	.addr_bytes_xip_0(\xip_controller|addr_bytes_xip[0]~0_combout ),
	.out_payload_0(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[0]~q ),
	.cmd_data_0(\xip_controller|cmd_data[0]~36_combout ),
	.mem_addr_reg_10(\xip_controller|mem_addr_reg[10]~q ),
	.mem_addr_reg_18(\xip_controller|mem_addr_reg[18]~q ),
	.mem_addr_reg_2(\xip_controller|mem_addr_reg[2]~q ),
	.out_payload_4(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[4]~q ),
	.cmd_data_4(\xip_controller|cmd_data[4]~43_combout ),
	.mem_addr_reg_8(\xip_controller|mem_addr_reg[8]~q ),
	.mem_addr_reg_16(\xip_controller|mem_addr_reg[16]~q ),
	.mem_addr_reg_0(\xip_controller|mem_addr_reg[0]~q ),
	.out_payload_2(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[2]~q ),
	.cmd_data_2(\xip_controller|cmd_data[2]~50_combout ),
	.mem_addr_reg_15(\xip_controller|mem_addr_reg[15]~q ),
	.mem_addr_reg_7(\xip_controller|mem_addr_reg[7]~q ),
	.WideOr19(\xip_controller|WideOr19~0_combout ),
	.out_payload_1(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[1]~q ),
	.cmd_data_1(\xip_controller|cmd_data[1]~57_combout ),
	.mem_addr_reg_17(\xip_controller|mem_addr_reg[17]~q ),
	.mem_addr_reg_9(\xip_controller|mem_addr_reg[9]~q ),
	.mem_addr_reg_1(\xip_controller|mem_addr_reg[1]~q ),
	.out_payload_3(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[3]~q ),
	.cmd_data_3(\xip_controller|cmd_data[3]~64_combout ),
	.mem_addr_reg_19(\xip_controller|mem_addr_reg[19]~q ),
	.mem_addr_reg_11(\xip_controller|mem_addr_reg[11]~q ),
	.mem_addr_reg_3(\xip_controller|mem_addr_reg[3]~q ),
	.out_payload_5(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[5]~q ),
	.cmd_data_5(\xip_controller|cmd_data[5]~71_combout ),
	.mem_addr_reg_12(\xip_controller|mem_addr_reg[12]~q ),
	.mem_addr_reg_20(\xip_controller|mem_addr_reg[20]~q ),
	.mem_addr_reg_4(\xip_controller|mem_addr_reg[4]~q ),
	.out_payload_6(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[6]~q ),
	.cmd_data_6(\xip_controller|cmd_data[6]~78_combout ),
	.mem_addr_reg_13(\xip_controller|mem_addr_reg[13]~q ),
	.mem_addr_reg_5(\xip_controller|mem_addr_reg[5]~q ),
	.out_payload_7(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[7]~q ),
	.cmd_data_7(\xip_controller|cmd_data[7]~85_combout ),
	.cmd_data_12(\xip_controller|cmd_data[12]~combout ),
	.out_payload_31(\xip_controller|avst_fifo_inst|avst_fifo|out_payload[31]~q ),
	.clk_clk(clk_clk),
	.avl_mem_read(avl_mem_read),
	.mem_burstcount({avl_mem_burstcount_6,avl_mem_burstcount_5,avl_mem_burstcount_4,avl_mem_burstcount_3,avl_mem_burstcount_2,avl_mem_burstcount_1,avl_mem_burstcount_0}),
	.avl_mem_write(avl_mem_write),
	.avl_mem_byteenable_0(avl_mem_byteenable_0),
	.avl_mem_byteenable_1(avl_mem_byteenable_1),
	.avl_mem_byteenable_2(avl_mem_byteenable_2),
	.avl_mem_byteenable_3(avl_mem_byteenable_3),
	.avl_mem_writedata_30(avl_mem_writedata_30),
	.avl_mem_writedata_29(avl_mem_writedata_29),
	.avl_mem_writedata_28(avl_mem_writedata_28),
	.avl_mem_writedata_27(avl_mem_writedata_27),
	.avl_mem_writedata_11(avl_mem_writedata_11),
	.avl_mem_writedata_18(avl_mem_writedata_18),
	.avl_mem_writedata_19(avl_mem_writedata_19),
	.avl_mem_writedata_21(avl_mem_writedata_21),
	.avl_mem_writedata_20(avl_mem_writedata_20),
	.avl_mem_writedata_22(avl_mem_writedata_22),
	.avl_mem_writedata_23(avl_mem_writedata_23),
	.avl_mem_writedata_24(avl_mem_writedata_24),
	.avl_mem_writedata_25(avl_mem_writedata_25),
	.avl_mem_writedata_26(avl_mem_writedata_26),
	.avl_mem_writedata_10(avl_mem_writedata_10),
	.avl_mem_writedata_8(avl_mem_writedata_8),
	.avl_mem_writedata_13(avl_mem_writedata_13),
	.avl_mem_writedata_17(avl_mem_writedata_17),
	.avl_mem_writedata_16(avl_mem_writedata_16),
	.avl_mem_writedata_15(avl_mem_writedata_15),
	.avl_mem_writedata_31(avl_mem_writedata_31),
	.avl_mem_writedata_14(avl_mem_writedata_14),
	.avl_mem_writedata_9(avl_mem_writedata_9),
	.mem_addr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_address_20,avl_mem_address_19,avl_mem_address_18,avl_mem_address_17,avl_mem_address_16,avl_mem_address_15,avl_mem_address_14,avl_mem_address_13,avl_mem_address_12,avl_mem_address_11,avl_mem_address_10,avl_mem_address_9,
avl_mem_address_8,avl_mem_address_7,avl_mem_address_6,avl_mem_address_5,avl_mem_address_4,avl_mem_address_3,avl_mem_address_2,avl_mem_address_1,avl_mem_address_0}),
	.avl_mem_writedata_0(avl_mem_writedata_0),
	.avl_mem_writedata_4(avl_mem_writedata_4),
	.avl_mem_writedata_12(avl_mem_writedata_12),
	.avl_mem_writedata_2(avl_mem_writedata_2),
	.avl_mem_writedata_1(avl_mem_writedata_1),
	.avl_mem_writedata_3(avl_mem_writedata_3),
	.avl_mem_writedata_5(avl_mem_writedata_5),
	.avl_mem_writedata_6(avl_mem_writedata_6),
	.avl_mem_writedata_7(avl_mem_writedata_7));

flashLoader_intel_generic_serial_flash_interface_csr csr_controller(
	.avl_rddata_local_0(avl_rddata_local_0),
	.avl_rddata_local_1(avl_rddata_local_1),
	.avl_rddata_local_2(avl_rddata_local_2),
	.avl_rddata_local_3(avl_rddata_local_3),
	.avl_rddata_local_4(avl_rddata_local_4),
	.avl_rddata_local_5(avl_rddata_local_5),
	.avl_rddata_local_6(avl_rddata_local_6),
	.avl_rddata_local_7(avl_rddata_local_7),
	.avl_rddata_local_8(avl_rddata_local_8),
	.avl_rddata_local_9(avl_rddata_local_9),
	.avl_rddata_local_10(avl_rddata_local_10),
	.avl_rddata_local_11(avl_rddata_local_11),
	.avl_rddata_local_12(avl_rddata_local_12),
	.avl_rddata_local_13(avl_rddata_local_13),
	.avl_rddata_local_14(avl_rddata_local_14),
	.avl_rddata_local_15(avl_rddata_local_15),
	.avl_rddata_local_16(avl_rddata_local_16),
	.avl_rddata_local_17(avl_rddata_local_17),
	.avl_rddata_local_18(avl_rddata_local_18),
	.avl_rddata_local_19(avl_rddata_local_19),
	.avl_rddata_local_20(avl_rddata_local_20),
	.avl_rddata_local_21(avl_rddata_local_21),
	.avl_rddata_local_22(avl_rddata_local_22),
	.avl_rddata_local_23(avl_rddata_local_23),
	.avl_rddata_local_24(avl_rddata_local_24),
	.avl_rddata_local_25(avl_rddata_local_25),
	.avl_rddata_local_26(avl_rddata_local_26),
	.avl_rddata_local_27(avl_rddata_local_27),
	.avl_rddata_local_28(avl_rddata_local_28),
	.avl_rddata_local_29(avl_rddata_local_29),
	.avl_rddata_local_30(avl_rddata_local_30),
	.avl_rddata_local_31(avl_rddata_local_31),
	.stateST_IDLE(\csr_controller|state.ST_IDLE~q ),
	.hold_waitrequest(\xip_controller|hold_waitrequest~q ),
	.csr_waitrequest1(csr_waitrequest),
	.avl_rddatavalid_local1(avl_rddatavalid_local),
	.csr_wr_inst_data_0(\csr_controller|csr_wr_inst_data[0]~q ),
	.csr_rd_inst_data_0(\csr_controller|csr_rd_inst_data[0]~q ),
	.csr_op_protocol_data_0(\csr_controller|csr_op_protocol_data[0]~q ),
	.csr_flash_cmd_wr_data_0_data_0(\csr_controller|csr_flash_cmd_wr_data_0_data[0]~q ),
	.csr_flash_cmd_addr_data_0(\csr_controller|csr_flash_cmd_addr_data[0]~q ),
	.csr_flash_cmd_wr_data_1_data_0(\csr_controller|csr_flash_cmd_wr_data_1_data[0]~q ),
	.csr_delay_setting_data_0(\csr_controller|csr_delay_setting_data[0]~q ),
	.csr_clk_baud_rate_data_0(\csr_controller|csr_clk_baud_rate_data[0]~q ),
	.csr_control_data_0(\csr_controller|csr_control_data[0]~q ),
	.csr_rd_capturing_data_0(\csr_controller|csr_rd_capturing_data[0]~q ),
	.reset(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.csr_wr_inst_data_1(\csr_controller|csr_wr_inst_data[1]~q ),
	.csr_rd_inst_data_1(\csr_controller|csr_rd_inst_data[1]~q ),
	.csr_op_protocol_data_1(\csr_controller|csr_op_protocol_data[1]~q ),
	.csr_flash_cmd_wr_data_0_data_1(\csr_controller|csr_flash_cmd_wr_data_0_data[1]~q ),
	.csr_flash_cmd_addr_data_1(\csr_controller|csr_flash_cmd_addr_data[1]~q ),
	.csr_flash_cmd_wr_data_1_data_1(\csr_controller|csr_flash_cmd_wr_data_1_data[1]~q ),
	.csr_delay_setting_data_1(\csr_controller|csr_delay_setting_data[1]~q ),
	.csr_clk_baud_rate_data_1(\csr_controller|csr_clk_baud_rate_data[1]~q ),
	.csr_rd_capturing_data_1(\csr_controller|csr_rd_capturing_data[1]~q ),
	.csr_wr_inst_data_2(\csr_controller|csr_wr_inst_data[2]~q ),
	.csr_rd_inst_data_2(\csr_controller|csr_rd_inst_data[2]~q ),
	.csr_flash_cmd_wr_data_0_data_2(\csr_controller|csr_flash_cmd_wr_data_0_data[2]~q ),
	.csr_flash_cmd_addr_data_2(\csr_controller|csr_flash_cmd_addr_data[2]~q ),
	.csr_flash_cmd_wr_data_1_data_2(\csr_controller|csr_flash_cmd_wr_data_1_data[2]~q ),
	.csr_delay_setting_data_2(\csr_controller|csr_delay_setting_data[2]~q ),
	.csr_clk_baud_rate_data_2(\csr_controller|csr_clk_baud_rate_data[2]~q ),
	.csr_rd_capturing_data_2(\csr_controller|csr_rd_capturing_data[2]~q ),
	.csr_wr_inst_data_3(\csr_controller|csr_wr_inst_data[3]~q ),
	.csr_rd_inst_data_3(\csr_controller|csr_rd_inst_data[3]~q ),
	.csr_flash_cmd_wr_data_0_data_3(\csr_controller|csr_flash_cmd_wr_data_0_data[3]~q ),
	.csr_flash_cmd_addr_data_3(\csr_controller|csr_flash_cmd_addr_data[3]~q ),
	.csr_flash_cmd_wr_data_1_data_3(\csr_controller|csr_flash_cmd_wr_data_1_data[3]~q ),
	.csr_delay_setting_data_3(\csr_controller|csr_delay_setting_data[3]~q ),
	.csr_clk_baud_rate_data_3(\csr_controller|csr_clk_baud_rate_data[3]~q ),
	.csr_rd_capturing_data_3(\csr_controller|csr_rd_capturing_data[3]~q ),
	.csr_wr_inst_data_4(\csr_controller|csr_wr_inst_data[4]~q ),
	.csr_delay_setting_data_4(\csr_controller|csr_delay_setting_data[4]~q ),
	.csr_flash_cmd_addr_data_4(\csr_controller|csr_flash_cmd_addr_data[4]~q ),
	.csr_op_protocol_data_4(\csr_controller|csr_op_protocol_data[4]~q ),
	.csr_clk_baud_rate_data_4(\csr_controller|csr_clk_baud_rate_data[4]~q ),
	.csr_control_data_4(\csr_controller|csr_control_data[4]~q ),
	.csr_rd_inst_data_4(\csr_controller|csr_rd_inst_data[4]~q ),
	.csr_flash_cmd_wr_data_1_data_4(\csr_controller|csr_flash_cmd_wr_data_1_data[4]~q ),
	.csr_flash_cmd_wr_data_0_data_4(\csr_controller|csr_flash_cmd_wr_data_0_data[4]~q ),
	.csr_delay_setting_data_5(\csr_controller|csr_delay_setting_data[5]~q ),
	.csr_wr_inst_data_5(\csr_controller|csr_wr_inst_data[5]~q ),
	.csr_rd_inst_data_5(\csr_controller|csr_rd_inst_data[5]~q ),
	.csr_op_protocol_data_5(\csr_controller|csr_op_protocol_data[5]~q ),
	.csr_control_data_5(\csr_controller|csr_control_data[5]~q ),
	.csr_flash_cmd_wr_data_1_data_5(\csr_controller|csr_flash_cmd_wr_data_1_data[5]~q ),
	.csr_flash_cmd_wr_data_0_data_5(\csr_controller|csr_flash_cmd_wr_data_0_data[5]~q ),
	.csr_flash_cmd_addr_data_5(\csr_controller|csr_flash_cmd_addr_data[5]~q ),
	.csr_wr_inst_data_6(\csr_controller|csr_wr_inst_data[6]~q ),
	.csr_rd_inst_data_6(\csr_controller|csr_rd_inst_data[6]~q ),
	.csr_delay_setting_data_6(\csr_controller|csr_delay_setting_data[6]~q ),
	.csr_control_data_6(\csr_controller|csr_control_data[6]~q ),
	.csr_flash_cmd_wr_data_1_data_6(\csr_controller|csr_flash_cmd_wr_data_1_data[6]~q ),
	.csr_flash_cmd_wr_data_0_data_6(\csr_controller|csr_flash_cmd_wr_data_0_data[6]~q ),
	.csr_flash_cmd_addr_data_6(\csr_controller|csr_flash_cmd_addr_data[6]~q ),
	.csr_delay_setting_data_7(\csr_controller|csr_delay_setting_data[7]~q ),
	.csr_wr_inst_data_7(\csr_controller|csr_wr_inst_data[7]~q ),
	.csr_rd_inst_data_7(\csr_controller|csr_rd_inst_data[7]~q ),
	.csr_control_data_7(\csr_controller|csr_control_data[7]~q ),
	.csr_flash_cmd_wr_data_1_data_7(\csr_controller|csr_flash_cmd_wr_data_1_data[7]~q ),
	.csr_flash_cmd_wr_data_0_data_7(\csr_controller|csr_flash_cmd_wr_data_0_data[7]~q ),
	.csr_flash_cmd_addr_data_7(\csr_controller|csr_flash_cmd_addr_data[7]~q ),
	.csr_rd_inst_data_8(\csr_controller|csr_rd_inst_data[8]~q ),
	.csr_op_protocol_data_8(\csr_controller|csr_op_protocol_data[8]~q ),
	.csr_flash_cmd_addr_data_8(\csr_controller|csr_flash_cmd_addr_data[8]~q ),
	.csr_control_data_8(\csr_controller|csr_control_data[8]~q ),
	.csr_flash_cmd_wr_data_0_data_8(\csr_controller|csr_flash_cmd_wr_data_0_data[8]~q ),
	.csr_wr_inst_data_8(\csr_controller|csr_wr_inst_data[8]~q ),
	.csr_flash_cmd_wr_data_1_data_8(\csr_controller|csr_flash_cmd_wr_data_1_data[8]~q ),
	.csr_flash_cmd_addr_data_9(\csr_controller|csr_flash_cmd_addr_data[9]~q ),
	.csr_rd_inst_data_9(\csr_controller|csr_rd_inst_data[9]~q ),
	.csr_op_protocol_data_9(\csr_controller|csr_op_protocol_data[9]~q ),
	.csr_flash_cmd_wr_data_0_data_9(\csr_controller|csr_flash_cmd_wr_data_0_data[9]~q ),
	.csr_wr_inst_data_9(\csr_controller|csr_wr_inst_data[9]~q ),
	.csr_flash_cmd_wr_data_1_data_9(\csr_controller|csr_flash_cmd_wr_data_1_data[9]~q ),
	.csr_rd_inst_data_10(\csr_controller|csr_rd_inst_data[10]~q ),
	.csr_flash_cmd_addr_data_10(\csr_controller|csr_flash_cmd_addr_data[10]~q ),
	.csr_flash_cmd_wr_data_0_data_10(\csr_controller|csr_flash_cmd_wr_data_0_data[10]~q ),
	.csr_wr_inst_data_10(\csr_controller|csr_wr_inst_data[10]~q ),
	.csr_flash_cmd_wr_data_1_data_10(\csr_controller|csr_flash_cmd_wr_data_1_data[10]~q ),
	.csr_flash_cmd_addr_data_11(\csr_controller|csr_flash_cmd_addr_data[11]~q ),
	.csr_rd_inst_data_11(\csr_controller|csr_rd_inst_data[11]~q ),
	.csr_flash_cmd_wr_data_0_data_11(\csr_controller|csr_flash_cmd_wr_data_0_data[11]~q ),
	.csr_wr_inst_data_11(\csr_controller|csr_wr_inst_data[11]~q ),
	.csr_flash_cmd_wr_data_1_data_11(\csr_controller|csr_flash_cmd_wr_data_1_data[11]~q ),
	.csr_rd_inst_data_12(\csr_controller|csr_rd_inst_data[12]~q ),
	.csr_op_protocol_data_12(\csr_controller|csr_op_protocol_data[12]~q ),
	.csr_flash_cmd_addr_data_12(\csr_controller|csr_flash_cmd_addr_data[12]~q ),
	.csr_flash_cmd_wr_data_0_data_12(\csr_controller|csr_flash_cmd_wr_data_0_data[12]~q ),
	.csr_wr_inst_data_12(\csr_controller|csr_wr_inst_data[12]~q ),
	.csr_flash_cmd_wr_data_1_data_12(\csr_controller|csr_flash_cmd_wr_data_1_data[12]~q ),
	.csr_flash_cmd_addr_data_13(\csr_controller|csr_flash_cmd_addr_data[13]~q ),
	.csr_op_protocol_data_13(\csr_controller|csr_op_protocol_data[13]~q ),
	.csr_flash_cmd_wr_data_0_data_13(\csr_controller|csr_flash_cmd_wr_data_0_data[13]~q ),
	.csr_wr_inst_data_13(\csr_controller|csr_wr_inst_data[13]~q ),
	.csr_flash_cmd_wr_data_1_data_13(\csr_controller|csr_flash_cmd_wr_data_1_data[13]~q ),
	.csr_flash_cmd_addr_data_14(\csr_controller|csr_flash_cmd_addr_data[14]~q ),
	.csr_flash_cmd_wr_data_0_data_14(\csr_controller|csr_flash_cmd_wr_data_0_data[14]~q ),
	.csr_wr_inst_data_14(\csr_controller|csr_wr_inst_data[14]~q ),
	.csr_flash_cmd_wr_data_1_data_14(\csr_controller|csr_flash_cmd_wr_data_1_data[14]~q ),
	.csr_flash_cmd_addr_data_15(\csr_controller|csr_flash_cmd_addr_data[15]~q ),
	.csr_flash_cmd_wr_data_0_data_15(\csr_controller|csr_flash_cmd_wr_data_0_data[15]~q ),
	.csr_wr_inst_data_15(\csr_controller|csr_wr_inst_data[15]~q ),
	.csr_flash_cmd_wr_data_1_data_15(\csr_controller|csr_flash_cmd_wr_data_1_data[15]~q ),
	.csr_op_protocol_data_16(\csr_controller|csr_op_protocol_data[16]~q ),
	.csr_flash_cmd_addr_data_16(\csr_controller|csr_flash_cmd_addr_data[16]~q ),
	.csr_flash_cmd_wr_data_0_data_16(\csr_controller|csr_flash_cmd_wr_data_0_data[16]~q ),
	.csr_flash_cmd_wr_data_1_data_16(\csr_controller|csr_flash_cmd_wr_data_1_data[16]~q ),
	.csr_flash_cmd_addr_data_17(\csr_controller|csr_flash_cmd_addr_data[17]~q ),
	.csr_op_protocol_data_17(\csr_controller|csr_op_protocol_data[17]~q ),
	.csr_flash_cmd_wr_data_0_data_17(\csr_controller|csr_flash_cmd_wr_data_0_data[17]~q ),
	.csr_flash_cmd_wr_data_1_data_17(\csr_controller|csr_flash_cmd_wr_data_1_data[17]~q ),
	.csr_flash_cmd_addr_data_18(\csr_controller|csr_flash_cmd_addr_data[18]~q ),
	.csr_flash_cmd_wr_data_0_data_18(\csr_controller|csr_flash_cmd_wr_data_0_data[18]~q ),
	.csr_flash_cmd_wr_data_1_data_18(\csr_controller|csr_flash_cmd_wr_data_1_data[18]~q ),
	.csr_flash_cmd_addr_data_19(\csr_controller|csr_flash_cmd_addr_data[19]~q ),
	.csr_flash_cmd_wr_data_0_data_19(\csr_controller|csr_flash_cmd_wr_data_0_data[19]~q ),
	.csr_flash_cmd_wr_data_1_data_19(\csr_controller|csr_flash_cmd_wr_data_1_data[19]~q ),
	.csr_flash_cmd_addr_data_20(\csr_controller|csr_flash_cmd_addr_data[20]~q ),
	.csr_flash_cmd_wr_data_0_data_20(\csr_controller|csr_flash_cmd_wr_data_0_data[20]~q ),
	.csr_flash_cmd_wr_data_1_data_20(\csr_controller|csr_flash_cmd_wr_data_1_data[20]~q ),
	.csr_flash_cmd_addr_data_21(\csr_controller|csr_flash_cmd_addr_data[21]~q ),
	.csr_flash_cmd_wr_data_0_data_21(\csr_controller|csr_flash_cmd_wr_data_0_data[21]~q ),
	.csr_flash_cmd_wr_data_1_data_21(\csr_controller|csr_flash_cmd_wr_data_1_data[21]~q ),
	.csr_flash_cmd_addr_data_22(\csr_controller|csr_flash_cmd_addr_data[22]~q ),
	.csr_flash_cmd_wr_data_0_data_22(\csr_controller|csr_flash_cmd_wr_data_0_data[22]~q ),
	.csr_flash_cmd_wr_data_1_data_22(\csr_controller|csr_flash_cmd_wr_data_1_data[22]~q ),
	.csr_flash_cmd_addr_data_23(\csr_controller|csr_flash_cmd_addr_data[23]~q ),
	.csr_flash_cmd_wr_data_0_data_23(\csr_controller|csr_flash_cmd_wr_data_0_data[23]~q ),
	.csr_flash_cmd_wr_data_1_data_23(\csr_controller|csr_flash_cmd_wr_data_1_data[23]~q ),
	.csr_flash_cmd_addr_data_24(\csr_controller|csr_flash_cmd_addr_data[24]~q ),
	.csr_flash_cmd_wr_data_0_data_24(\csr_controller|csr_flash_cmd_wr_data_0_data[24]~q ),
	.csr_flash_cmd_wr_data_1_data_24(\csr_controller|csr_flash_cmd_wr_data_1_data[24]~q ),
	.csr_flash_cmd_addr_data_25(\csr_controller|csr_flash_cmd_addr_data[25]~q ),
	.csr_flash_cmd_wr_data_0_data_25(\csr_controller|csr_flash_cmd_wr_data_0_data[25]~q ),
	.csr_flash_cmd_wr_data_1_data_25(\csr_controller|csr_flash_cmd_wr_data_1_data[25]~q ),
	.csr_flash_cmd_addr_data_26(\csr_controller|csr_flash_cmd_addr_data[26]~q ),
	.csr_flash_cmd_wr_data_0_data_26(\csr_controller|csr_flash_cmd_wr_data_0_data[26]~q ),
	.csr_flash_cmd_wr_data_1_data_26(\csr_controller|csr_flash_cmd_wr_data_1_data[26]~q ),
	.csr_flash_cmd_addr_data_27(\csr_controller|csr_flash_cmd_addr_data[27]~q ),
	.csr_flash_cmd_wr_data_0_data_27(\csr_controller|csr_flash_cmd_wr_data_0_data[27]~q ),
	.csr_flash_cmd_wr_data_1_data_27(\csr_controller|csr_flash_cmd_wr_data_1_data[27]~q ),
	.csr_flash_cmd_addr_data_28(\csr_controller|csr_flash_cmd_addr_data[28]~q ),
	.csr_flash_cmd_wr_data_0_data_28(\csr_controller|csr_flash_cmd_wr_data_0_data[28]~q ),
	.csr_flash_cmd_wr_data_1_data_28(\csr_controller|csr_flash_cmd_wr_data_1_data[28]~q ),
	.csr_flash_cmd_addr_data_29(\csr_controller|csr_flash_cmd_addr_data[29]~q ),
	.csr_flash_cmd_wr_data_0_data_29(\csr_controller|csr_flash_cmd_wr_data_0_data[29]~q ),
	.csr_flash_cmd_wr_data_1_data_29(\csr_controller|csr_flash_cmd_wr_data_1_data[29]~q ),
	.csr_flash_cmd_addr_data_30(\csr_controller|csr_flash_cmd_addr_data[30]~q ),
	.csr_flash_cmd_wr_data_0_data_30(\csr_controller|csr_flash_cmd_wr_data_0_data[30]~q ),
	.csr_flash_cmd_wr_data_1_data_30(\csr_controller|csr_flash_cmd_wr_data_1_data[30]~q ),
	.csr_flash_cmd_addr_data_31(\csr_controller|csr_flash_cmd_addr_data[31]~q ),
	.csr_flash_cmd_wr_data_0_data_31(\csr_controller|csr_flash_cmd_wr_data_0_data[31]~q ),
	.csr_flash_cmd_wr_data_1_data_31(\csr_controller|csr_flash_cmd_wr_data_1_data[31]~q ),
	.stateST_SEND_DUMMY_RSP(\serial_flash_inf_cmd_gen_inst|state.ST_SEND_DUMMY_RSP~q ),
	.out_valid(\serial_flash_inf_cmd_gen_inst|data_adapter_8_32_inst|out_valid~q ),
	.out_endofpacket(\serial_flash_inf_cmd_gen_inst|data_adapter_8_32_inst|out_endofpacket~q ),
	.in_cmd_channel_reg_1(\serial_flash_inf_cmd_gen_inst|in_cmd_channel_reg[1]~q ),
	.stateST_WAIT_RSP(\csr_controller|state.ST_WAIT_RSP~q ),
	.sink_ready(\merlin_demultiplexer_0|sink_ready~0_combout ),
	.out_rsp_data_0(\serial_flash_inf_cmd_gen_inst|out_rsp_data[0]~0_combout ),
	.out_rsp_data_1(\serial_flash_inf_cmd_gen_inst|out_rsp_data[1]~1_combout ),
	.out_rsp_data_2(\serial_flash_inf_cmd_gen_inst|out_rsp_data[2]~2_combout ),
	.out_rsp_data_3(\serial_flash_inf_cmd_gen_inst|out_rsp_data[3]~3_combout ),
	.out_rsp_data_4(\serial_flash_inf_cmd_gen_inst|out_rsp_data[4]~4_combout ),
	.out_rsp_data_5(\serial_flash_inf_cmd_gen_inst|out_rsp_data[5]~5_combout ),
	.out_rsp_data_6(\serial_flash_inf_cmd_gen_inst|out_rsp_data[6]~6_combout ),
	.out_rsp_data_7(\serial_flash_inf_cmd_gen_inst|out_rsp_data[7]~7_combout ),
	.out_rsp_data_8(\serial_flash_inf_cmd_gen_inst|out_rsp_data[8]~8_combout ),
	.out_rsp_data_9(\serial_flash_inf_cmd_gen_inst|out_rsp_data[9]~9_combout ),
	.out_rsp_data_10(\serial_flash_inf_cmd_gen_inst|out_rsp_data[10]~10_combout ),
	.out_rsp_data_11(\serial_flash_inf_cmd_gen_inst|out_rsp_data[11]~11_combout ),
	.out_rsp_data_12(\serial_flash_inf_cmd_gen_inst|out_rsp_data[12]~12_combout ),
	.out_rsp_data_13(\serial_flash_inf_cmd_gen_inst|out_rsp_data[13]~13_combout ),
	.out_rsp_data_14(\serial_flash_inf_cmd_gen_inst|out_rsp_data[14]~14_combout ),
	.out_rsp_data_15(\serial_flash_inf_cmd_gen_inst|out_rsp_data[15]~15_combout ),
	.out_rsp_data_16(\serial_flash_inf_cmd_gen_inst|out_rsp_data[16]~16_combout ),
	.out_rsp_data_17(\serial_flash_inf_cmd_gen_inst|out_rsp_data[17]~17_combout ),
	.out_rsp_data_18(\serial_flash_inf_cmd_gen_inst|out_rsp_data[18]~18_combout ),
	.out_rsp_data_19(\serial_flash_inf_cmd_gen_inst|out_rsp_data[19]~19_combout ),
	.out_rsp_data_20(\serial_flash_inf_cmd_gen_inst|out_rsp_data[20]~20_combout ),
	.out_rsp_data_21(\serial_flash_inf_cmd_gen_inst|out_rsp_data[21]~21_combout ),
	.out_rsp_data_22(\serial_flash_inf_cmd_gen_inst|out_rsp_data[22]~22_combout ),
	.out_rsp_data_23(\serial_flash_inf_cmd_gen_inst|out_rsp_data[23]~23_combout ),
	.out_rsp_data_24(\serial_flash_inf_cmd_gen_inst|out_rsp_data[24]~24_combout ),
	.out_rsp_data_25(\serial_flash_inf_cmd_gen_inst|out_rsp_data[25]~25_combout ),
	.out_rsp_data_26(\serial_flash_inf_cmd_gen_inst|out_rsp_data[26]~26_combout ),
	.out_rsp_data_27(\serial_flash_inf_cmd_gen_inst|out_rsp_data[27]~27_combout ),
	.out_rsp_data_28(\serial_flash_inf_cmd_gen_inst|out_rsp_data[28]~28_combout ),
	.out_rsp_data_29(\serial_flash_inf_cmd_gen_inst|out_rsp_data[29]~29_combout ),
	.out_rsp_data_30(\serial_flash_inf_cmd_gen_inst|out_rsp_data[30]~30_combout ),
	.out_rsp_data_31(\serial_flash_inf_cmd_gen_inst|out_rsp_data[31]~31_combout ),
	.saved_grant_1(\multiplexer|saved_grant[1]~q ),
	.stateST_SEND_HEADER(\csr_controller|state.ST_SEND_HEADER~q ),
	.stateST_SEND_DATA_1(\csr_controller|state.ST_SEND_DATA_1~q ),
	.stateST_SEND_DATA_0(\csr_controller|state.ST_SEND_DATA_0~q ),
	.has_data_in1(\csr_controller|has_data_in~q ),
	.more_than_4bytes_data1(\csr_controller|more_than_4bytes_data~q ),
	.src_payload_0(\multiplexer|src_payload[0]~1_combout ),
	.Selector18(\serial_flash_inf_cmd_gen_inst|Selector18~5_combout ),
	.sink1_ready(\multiplexer|sink1_ready~combout ),
	.Selector34(\csr_controller|Selector34~0_combout ),
	.has_data_out1(\csr_controller|has_data_out~q ),
	.numb_data_0(\csr_controller|numb_data[0]~q ),
	.numb_data_1(\csr_controller|numb_data[1]~q ),
	.numb_data_3(\csr_controller|numb_data[3]~q ),
	.numb_data_2(\csr_controller|numb_data[2]~q ),
	.has_addr1(\csr_controller|has_addr~q ),
	.numb_dummy_0(\csr_controller|numb_dummy[0]~q ),
	.numb_dummy_4(\csr_controller|numb_dummy[4]~q ),
	.numb_dummy_3(\csr_controller|numb_dummy[3]~q ),
	.numb_dummy_2(\csr_controller|numb_dummy[2]~q ),
	.numb_dummy_1(\csr_controller|numb_dummy[1]~q ),
	.is_4bytes_addr1(\csr_controller|is_4bytes_addr~q ),
	.opcode_0(\csr_controller|opcode[0]~q ),
	.opcode_4(\csr_controller|opcode[4]~q ),
	.opcode_2(\csr_controller|opcode[2]~q ),
	.opcode_1(\csr_controller|opcode[1]~q ),
	.opcode_3(\csr_controller|opcode[3]~q ),
	.opcode_5(\csr_controller|opcode[5]~q ),
	.opcode_6(\csr_controller|opcode[6]~q ),
	.opcode_7(\csr_controller|opcode[7]~q ),
	.has_dummy1(\csr_controller|has_dummy~q ),
	.avl_csr_address_1(avl_csr_address_1),
	.avl_csr_address_0(avl_csr_address_0),
	.avl_csr_address_2(avl_csr_address_2),
	.avl_csr_address_3(avl_csr_address_3),
	.avl_csr_read(avl_csr_read),
	.avl_csr_address_4(avl_csr_address_4),
	.avl_csr_address_5(avl_csr_address_5),
	.clk(clk_clk),
	.avl_csr_write(avl_csr_write),
	.csr_wrdata({avl_csr_writedata_31,avl_csr_writedata_30,avl_csr_writedata_29,avl_csr_writedata_28,avl_csr_writedata_27,avl_csr_writedata_26,avl_csr_writedata_25,avl_csr_writedata_24,avl_csr_writedata_23,avl_csr_writedata_22,avl_csr_writedata_21,avl_csr_writedata_20,
avl_csr_writedata_19,avl_csr_writedata_18,avl_csr_writedata_17,avl_csr_writedata_16,avl_csr_writedata_15,avl_csr_writedata_14,avl_csr_writedata_13,avl_csr_writedata_12,avl_csr_writedata_11,avl_csr_writedata_10,avl_csr_writedata_9,avl_csr_writedata_8,
avl_csr_writedata_7,avl_csr_writedata_6,avl_csr_writedata_5,avl_csr_writedata_4,avl_csr_writedata_3,avl_csr_writedata_2,avl_csr_writedata_1,avl_csr_writedata_0}));

endmodule

module flashLoader_altera_reset_controller (
	altera_reset_synchronizer_int_chain_out,
	clk_clk,
	reset_reset)/* synthesis synthesis_greybox=0 */;
output 	altera_reset_synchronizer_int_chain_out;
input 	clk_clk;
input 	reset_reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



flashLoader_altera_reset_synchronizer_1 alt_rst_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(altera_reset_synchronizer_int_chain_out),
	.clk(clk_clk),
	.reset_reset(reset_reset));

endmodule

module flashLoader_altera_reset_synchronizer_1 (
	altera_reset_synchronizer_int_chain_out1,
	clk,
	reset_reset)/* synthesis synthesis_greybox=0 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;
input 	reset_reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(!reset_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!reset_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(!reset_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module flashLoader_flashLoader_intel_generic_serial_flash_interface_top_0_merlin_demultiplexer_0 (
	in_cmd_channel_reg_1,
	stateST_WAIT_RSP,
	sink_ready,
	in_cmd_channel_reg_0,
	WideOr01)/* synthesis synthesis_greybox=0 */;
input 	in_cmd_channel_reg_1;
input 	stateST_WAIT_RSP;
output 	sink_ready;
input 	in_cmd_channel_reg_0;
output 	WideOr01;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \sink_ready~0 (
	.dataa(in_cmd_channel_reg_1),
	.datab(stateST_WAIT_RSP),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(sink_ready),
	.cout());
defparam \sink_ready~0 .lut_mask = 16'h8888;
defparam \sink_ready~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb WideOr0(
	.dataa(in_cmd_channel_reg_0),
	.datab(in_cmd_channel_reg_1),
	.datac(stateST_WAIT_RSP),
	.datad(gnd),
	.cin(gnd),
	.combout(WideOr01),
	.cout());
defparam WideOr0.lut_mask = 16'hEAEA;
defparam WideOr0.sum_lutc_input = "datac";

endmodule

module flashLoader_flashLoader_intel_generic_serial_flash_interface_top_0_multiplexer (
	stateST_IDLE,
	csr_flash_cmd_wr_data_0_data_0,
	csr_flash_cmd_wr_data_1_data_0,
	altera_reset_synchronizer_int_chain_out,
	csr_flash_cmd_wr_data_0_data_1,
	csr_flash_cmd_wr_data_1_data_1,
	csr_flash_cmd_wr_data_0_data_2,
	csr_flash_cmd_wr_data_1_data_2,
	csr_flash_cmd_wr_data_0_data_3,
	csr_flash_cmd_wr_data_1_data_3,
	csr_control_data_4,
	csr_flash_cmd_wr_data_1_data_4,
	csr_flash_cmd_wr_data_0_data_4,
	csr_control_data_5,
	csr_flash_cmd_wr_data_1_data_5,
	csr_flash_cmd_wr_data_0_data_5,
	csr_control_data_6,
	csr_flash_cmd_wr_data_1_data_6,
	csr_flash_cmd_wr_data_0_data_6,
	csr_control_data_7,
	csr_flash_cmd_wr_data_1_data_7,
	csr_flash_cmd_wr_data_0_data_7,
	csr_flash_cmd_wr_data_0_data_8,
	csr_flash_cmd_wr_data_1_data_8,
	csr_flash_cmd_wr_data_0_data_9,
	csr_flash_cmd_wr_data_1_data_9,
	csr_flash_cmd_wr_data_0_data_10,
	csr_flash_cmd_wr_data_1_data_10,
	csr_rd_inst_data_11,
	csr_flash_cmd_wr_data_0_data_11,
	csr_flash_cmd_wr_data_1_data_11,
	csr_rd_inst_data_12,
	csr_flash_cmd_wr_data_0_data_13,
	csr_flash_cmd_wr_data_1_data_13,
	csr_flash_cmd_wr_data_0_data_14,
	csr_flash_cmd_wr_data_1_data_14,
	csr_flash_cmd_wr_data_0_data_15,
	csr_flash_cmd_wr_data_1_data_15,
	csr_flash_cmd_wr_data_0_data_16,
	csr_flash_cmd_wr_data_1_data_16,
	csr_flash_cmd_wr_data_0_data_17,
	csr_flash_cmd_wr_data_1_data_17,
	csr_flash_cmd_wr_data_0_data_18,
	csr_flash_cmd_wr_data_1_data_18,
	csr_flash_cmd_wr_data_0_data_19,
	csr_flash_cmd_wr_data_1_data_19,
	csr_flash_cmd_wr_data_0_data_20,
	csr_flash_cmd_wr_data_1_data_20,
	csr_flash_cmd_wr_data_0_data_21,
	csr_flash_cmd_wr_data_1_data_21,
	csr_flash_cmd_wr_data_0_data_22,
	csr_flash_cmd_wr_data_1_data_22,
	csr_flash_cmd_wr_data_0_data_23,
	csr_flash_cmd_wr_data_1_data_23,
	csr_flash_cmd_wr_data_0_data_24,
	csr_flash_cmd_wr_data_1_data_24,
	csr_flash_cmd_wr_data_0_data_25,
	csr_flash_cmd_wr_data_1_data_25,
	csr_flash_cmd_wr_data_0_data_26,
	csr_flash_cmd_wr_data_1_data_26,
	csr_flash_cmd_wr_data_0_data_27,
	csr_flash_cmd_wr_data_1_data_27,
	csr_flash_cmd_wr_data_0_data_28,
	csr_flash_cmd_wr_data_1_data_28,
	csr_flash_cmd_wr_data_0_data_29,
	csr_flash_cmd_wr_data_1_data_29,
	csr_flash_cmd_wr_data_0_data_30,
	csr_flash_cmd_wr_data_1_data_30,
	stateST_WAIT_RSP,
	saved_grant_1,
	stateST_SEND_HEADER,
	saved_grant_0,
	current_stateSTATE_WR_CMD,
	current_stateSTATE_STATUS_CMD,
	current_stateSTATE_POLL_CMD,
	current_stateSTATE_READ_CMD,
	WideOr13,
	src_startofpacket1,
	src_valid,
	current_stateSTATE_WR_DATA,
	cmd_valid,
	stateST_SEND_DATA,
	Selector18,
	WideOr0,
	in_ready,
	WideOr01,
	adap_out_cmd_ready,
	Selector181,
	stateST_SEND_DATA_1,
	stateST_SEND_DATA_0,
	has_data_in,
	more_than_4bytes_data,
	src_payload_0,
	Selector182,
	sink0_ready,
	src_data_30,
	is_burst_reg,
	mem_write_data_reg_30,
	mem_byteenable_reg_0,
	mem_byteenable_reg_3,
	mem_byteenable_reg_2,
	mem_byteenable_reg_1,
	src_data_301,
	out_payload_30,
	cmd_valid1,
	src_data_302,
	src_data_303,
	src_data_29,
	mem_write_data_reg_29,
	out_payload_29,
	src_data_291,
	src_data_292,
	src_data_28,
	mem_write_data_reg_28,
	out_payload_28,
	src_data_281,
	src_data_282,
	src_data_27,
	mem_write_data_reg_27,
	out_payload_27,
	src_data_271,
	src_data_272,
	WideOr11,
	out_payload_32,
	src_payload_01,
	sink1_ready1,
	Selector34,
	has_data_out,
	src_data_11,
	cmd_data_11,
	src_data_111,
	numb_data_0,
	Add1,
	Selector20,
	out_payload_18,
	mem_write_data_reg_18,
	src_data_18,
	numb_data_1,
	src_data_19,
	Add11,
	mem_write_data_reg_19,
	out_payload_19,
	src_data_191,
	src_data_192,
	numb_data_3,
	src_data_21,
	mem_write_data_reg_21,
	out_payload_21,
	mem_burstcount_reg_1,
	src_data_211,
	src_data_212,
	numb_data_2,
	src_data_20,
	mem_write_data_reg_20,
	out_payload_20,
	mem_burstcount_reg_0,
	src_data_201,
	src_data_202,
	mem_write_data_reg_22,
	out_payload_22,
	mem_burstcount_reg_2,
	src_data_22,
	mem_write_data_reg_23,
	out_payload_23,
	mem_burstcount_reg_3,
	src_data_23,
	mem_write_data_reg_24,
	out_payload_24,
	mem_burstcount_reg_4,
	src_data_24,
	mem_write_data_reg_25,
	out_payload_25,
	mem_burstcount_reg_5,
	src_data_25,
	mem_write_data_reg_26,
	out_payload_26,
	mem_burstcount_reg_6,
	src_data_26,
	src_data_10,
	cmd_data_10,
	src_data_101,
	has_addr,
	src_data_8,
	cmd_data_8,
	src_data_81,
	numb_dummy_0,
	src_data_13,
	cmd_data_13,
	src_data_131,
	numb_dummy_4,
	src_data_17,
	mem_write_data_reg_17,
	out_payload_17,
	src_data_171,
	src_data_172,
	numb_dummy_3,
	src_data_16,
	mem_write_data_reg_16,
	out_payload_16,
	src_data_161,
	src_data_162,
	numb_dummy_2,
	src_data_15,
	cmd_data_15,
	src_data_151,
	numb_dummy_1,
	src_data_14,
	cmd_data_14,
	src_data_141,
	is_4bytes_addr,
	src_data_9,
	cmd_data_9,
	src_data_91,
	opcode_0,
	out_payload_0,
	cmd_data_0,
	src_data_0,
	opcode_4,
	out_payload_4,
	cmd_data_4,
	src_data_4,
	opcode_2,
	out_payload_2,
	cmd_data_2,
	src_data_2,
	opcode_1,
	out_payload_1,
	cmd_data_1,
	src_data_1,
	opcode_3,
	out_payload_3,
	cmd_data_3,
	src_data_3,
	opcode_5,
	out_payload_5,
	cmd_data_5,
	src_data_5,
	opcode_6,
	out_payload_6,
	cmd_data_6,
	src_data_6,
	opcode_7,
	out_payload_7,
	cmd_data_7,
	src_data_7,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	stateST_IDLE;
input 	csr_flash_cmd_wr_data_0_data_0;
input 	csr_flash_cmd_wr_data_1_data_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	csr_flash_cmd_wr_data_0_data_1;
input 	csr_flash_cmd_wr_data_1_data_1;
input 	csr_flash_cmd_wr_data_0_data_2;
input 	csr_flash_cmd_wr_data_1_data_2;
input 	csr_flash_cmd_wr_data_0_data_3;
input 	csr_flash_cmd_wr_data_1_data_3;
input 	csr_control_data_4;
input 	csr_flash_cmd_wr_data_1_data_4;
input 	csr_flash_cmd_wr_data_0_data_4;
input 	csr_control_data_5;
input 	csr_flash_cmd_wr_data_1_data_5;
input 	csr_flash_cmd_wr_data_0_data_5;
input 	csr_control_data_6;
input 	csr_flash_cmd_wr_data_1_data_6;
input 	csr_flash_cmd_wr_data_0_data_6;
input 	csr_control_data_7;
input 	csr_flash_cmd_wr_data_1_data_7;
input 	csr_flash_cmd_wr_data_0_data_7;
input 	csr_flash_cmd_wr_data_0_data_8;
input 	csr_flash_cmd_wr_data_1_data_8;
input 	csr_flash_cmd_wr_data_0_data_9;
input 	csr_flash_cmd_wr_data_1_data_9;
input 	csr_flash_cmd_wr_data_0_data_10;
input 	csr_flash_cmd_wr_data_1_data_10;
input 	csr_rd_inst_data_11;
input 	csr_flash_cmd_wr_data_0_data_11;
input 	csr_flash_cmd_wr_data_1_data_11;
input 	csr_rd_inst_data_12;
input 	csr_flash_cmd_wr_data_0_data_13;
input 	csr_flash_cmd_wr_data_1_data_13;
input 	csr_flash_cmd_wr_data_0_data_14;
input 	csr_flash_cmd_wr_data_1_data_14;
input 	csr_flash_cmd_wr_data_0_data_15;
input 	csr_flash_cmd_wr_data_1_data_15;
input 	csr_flash_cmd_wr_data_0_data_16;
input 	csr_flash_cmd_wr_data_1_data_16;
input 	csr_flash_cmd_wr_data_0_data_17;
input 	csr_flash_cmd_wr_data_1_data_17;
input 	csr_flash_cmd_wr_data_0_data_18;
input 	csr_flash_cmd_wr_data_1_data_18;
input 	csr_flash_cmd_wr_data_0_data_19;
input 	csr_flash_cmd_wr_data_1_data_19;
input 	csr_flash_cmd_wr_data_0_data_20;
input 	csr_flash_cmd_wr_data_1_data_20;
input 	csr_flash_cmd_wr_data_0_data_21;
input 	csr_flash_cmd_wr_data_1_data_21;
input 	csr_flash_cmd_wr_data_0_data_22;
input 	csr_flash_cmd_wr_data_1_data_22;
input 	csr_flash_cmd_wr_data_0_data_23;
input 	csr_flash_cmd_wr_data_1_data_23;
input 	csr_flash_cmd_wr_data_0_data_24;
input 	csr_flash_cmd_wr_data_1_data_24;
input 	csr_flash_cmd_wr_data_0_data_25;
input 	csr_flash_cmd_wr_data_1_data_25;
input 	csr_flash_cmd_wr_data_0_data_26;
input 	csr_flash_cmd_wr_data_1_data_26;
input 	csr_flash_cmd_wr_data_0_data_27;
input 	csr_flash_cmd_wr_data_1_data_27;
input 	csr_flash_cmd_wr_data_0_data_28;
input 	csr_flash_cmd_wr_data_1_data_28;
input 	csr_flash_cmd_wr_data_0_data_29;
input 	csr_flash_cmd_wr_data_1_data_29;
input 	csr_flash_cmd_wr_data_0_data_30;
input 	csr_flash_cmd_wr_data_1_data_30;
input 	stateST_WAIT_RSP;
output 	saved_grant_1;
input 	stateST_SEND_HEADER;
output 	saved_grant_0;
input 	current_stateSTATE_WR_CMD;
input 	current_stateSTATE_STATUS_CMD;
input 	current_stateSTATE_POLL_CMD;
input 	current_stateSTATE_READ_CMD;
input 	WideOr13;
output 	src_startofpacket1;
output 	src_valid;
input 	current_stateSTATE_WR_DATA;
input 	cmd_valid;
input 	stateST_SEND_DATA;
input 	Selector18;
input 	WideOr0;
input 	in_ready;
input 	WideOr01;
input 	adap_out_cmd_ready;
input 	Selector181;
input 	stateST_SEND_DATA_1;
input 	stateST_SEND_DATA_0;
input 	has_data_in;
input 	more_than_4bytes_data;
output 	src_payload_0;
input 	Selector182;
output 	sink0_ready;
output 	src_data_30;
input 	is_burst_reg;
input 	mem_write_data_reg_30;
input 	mem_byteenable_reg_0;
input 	mem_byteenable_reg_3;
input 	mem_byteenable_reg_2;
input 	mem_byteenable_reg_1;
output 	src_data_301;
input 	out_payload_30;
input 	cmd_valid1;
output 	src_data_302;
output 	src_data_303;
output 	src_data_29;
input 	mem_write_data_reg_29;
input 	out_payload_29;
output 	src_data_291;
output 	src_data_292;
output 	src_data_28;
input 	mem_write_data_reg_28;
input 	out_payload_28;
output 	src_data_281;
output 	src_data_282;
output 	src_data_27;
input 	mem_write_data_reg_27;
input 	out_payload_27;
output 	src_data_271;
output 	src_data_272;
output 	WideOr11;
input 	out_payload_32;
output 	src_payload_01;
output 	sink1_ready1;
input 	Selector34;
input 	has_data_out;
output 	src_data_11;
input 	cmd_data_11;
output 	src_data_111;
input 	numb_data_0;
input 	Add1;
input 	Selector20;
input 	out_payload_18;
input 	mem_write_data_reg_18;
output 	src_data_18;
input 	numb_data_1;
output 	src_data_19;
input 	Add11;
input 	mem_write_data_reg_19;
input 	out_payload_19;
output 	src_data_191;
output 	src_data_192;
input 	numb_data_3;
output 	src_data_21;
input 	mem_write_data_reg_21;
input 	out_payload_21;
input 	mem_burstcount_reg_1;
output 	src_data_211;
output 	src_data_212;
input 	numb_data_2;
output 	src_data_20;
input 	mem_write_data_reg_20;
input 	out_payload_20;
input 	mem_burstcount_reg_0;
output 	src_data_201;
output 	src_data_202;
input 	mem_write_data_reg_22;
input 	out_payload_22;
input 	mem_burstcount_reg_2;
output 	src_data_22;
input 	mem_write_data_reg_23;
input 	out_payload_23;
input 	mem_burstcount_reg_3;
output 	src_data_23;
input 	mem_write_data_reg_24;
input 	out_payload_24;
input 	mem_burstcount_reg_4;
output 	src_data_24;
input 	mem_write_data_reg_25;
input 	out_payload_25;
input 	mem_burstcount_reg_5;
output 	src_data_25;
input 	mem_write_data_reg_26;
input 	out_payload_26;
input 	mem_burstcount_reg_6;
output 	src_data_26;
output 	src_data_10;
input 	cmd_data_10;
output 	src_data_101;
input 	has_addr;
output 	src_data_8;
input 	cmd_data_8;
output 	src_data_81;
input 	numb_dummy_0;
output 	src_data_13;
input 	cmd_data_13;
output 	src_data_131;
input 	numb_dummy_4;
output 	src_data_17;
input 	mem_write_data_reg_17;
input 	out_payload_17;
output 	src_data_171;
output 	src_data_172;
input 	numb_dummy_3;
output 	src_data_16;
input 	mem_write_data_reg_16;
input 	out_payload_16;
output 	src_data_161;
output 	src_data_162;
input 	numb_dummy_2;
output 	src_data_15;
input 	cmd_data_15;
output 	src_data_151;
input 	numb_dummy_1;
output 	src_data_14;
input 	cmd_data_14;
output 	src_data_141;
input 	is_4bytes_addr;
output 	src_data_9;
input 	cmd_data_9;
output 	src_data_91;
input 	opcode_0;
input 	out_payload_0;
input 	cmd_data_0;
output 	src_data_0;
input 	opcode_4;
input 	out_payload_4;
input 	cmd_data_4;
output 	src_data_4;
input 	opcode_2;
input 	out_payload_2;
input 	cmd_data_2;
output 	src_data_2;
input 	opcode_1;
input 	out_payload_1;
input 	cmd_data_1;
output 	src_data_1;
input 	opcode_3;
input 	out_payload_3;
input 	cmd_data_3;
output 	src_data_3;
input 	opcode_5;
input 	out_payload_5;
input 	cmd_data_5;
output 	src_data_5;
input 	opcode_6;
input 	out_payload_6;
input 	cmd_data_6;
output 	src_data_6;
input 	opcode_7;
input 	out_payload_7;
input 	cmd_data_7;
output 	src_data_7;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[1]~0_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;
wire \src_payload~0_combout ;
wire \sink0_ready~0_combout ;
wire \src_data[30]~2_combout ;
wire \src_data[30]~4_combout ;
wire \src_data[30]~6_combout ;
wire \src_data[29]~9_combout ;
wire \src_data[29]~11_combout ;
wire \src_data[28]~14_combout ;
wire \src_data[28]~16_combout ;
wire \src_data[27]~19_combout ;
wire \src_data[27]~21_combout ;
wire \src_payload[0]~2_combout ;
wire \src_data[11]~24_combout ;
wire \src_data[18]~27_combout ;
wire \src_data[18]~28_combout ;
wire \src_data[18]~124_combout ;
wire \src_data[18]~29_combout ;
wire \src_data[18]~30_combout ;
wire \src_data[18]~31_combout ;
wire \src_data[19]~33_combout ;
wire \src_data[19]~35_combout ;
wire \src_data[19]~36_combout ;
wire \src_data[21]~39_combout ;
wire \src_data[21]~41_combout ;
wire \src_data[21]~42_combout ;
wire \src_data[20]~45_combout ;
wire \src_data[20]~47_combout ;
wire \src_data[20]~48_combout ;
wire \src_data[20]~49_combout ;
wire \src_data[22]~52_combout ;
wire \src_data[22]~53_combout ;
wire \src_data[22]~54_combout ;
wire \src_data[23]~56_combout ;
wire \src_data[23]~57_combout ;
wire \src_data[23]~58_combout ;
wire \src_data[24]~60_combout ;
wire \src_data[24]~61_combout ;
wire \src_data[24]~62_combout ;
wire \src_data[25]~64_combout ;
wire \src_data[25]~65_combout ;
wire \src_data[25]~66_combout ;
wire \src_data[26]~68_combout ;
wire \src_data[26]~69_combout ;
wire \src_data[26]~70_combout ;
wire \src_data[10]~72_combout ;
wire \src_data[8]~75_combout ;
wire \src_data[13]~78_combout ;
wire \src_data[17]~81_combout ;
wire \src_data[17]~83_combout ;
wire \src_data[16]~86_combout ;
wire \src_data[16]~88_combout ;
wire \src_data[15]~91_combout ;
wire \src_data[14]~94_combout ;
wire \src_data[9]~97_combout ;
wire \src_data[0]~100_combout ;
wire \src_data[0]~101_combout ;
wire \src_payload~4_combout ;
wire \src_payload~5_combout ;
wire \src_data[4]~103_combout ;
wire \src_data[4]~104_combout ;
wire \src_payload~6_combout ;
wire \src_data[2]~106_combout ;
wire \src_data[2]~107_combout ;
wire \src_payload~7_combout ;
wire \src_data[1]~109_combout ;
wire \src_data[1]~110_combout ;
wire \src_payload~8_combout ;
wire \src_data[3]~112_combout ;
wire \src_data[3]~113_combout ;
wire \src_payload~9_combout ;
wire \src_data[5]~115_combout ;
wire \src_data[5]~116_combout ;
wire \src_payload~10_combout ;
wire \src_data[6]~118_combout ;
wire \src_data[6]~119_combout ;
wire \src_payload~11_combout ;
wire \src_data[7]~121_combout ;
wire \src_data[7]~122_combout ;
wire \src_payload~12_combout ;


flashLoader_altera_merlin_arbitrator arb(
	.stateST_IDLE(stateST_IDLE),
	.stateST_WAIT_RSP(stateST_WAIT_RSP),
	.cmd_valid(cmd_valid),
	.grant_1(\arb|grant[1]~0_combout ));

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(cmd_valid),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

cycloneive_lcell_comb src_startofpacket(
	.dataa(\src_payload~0_combout ),
	.datab(saved_grant_0),
	.datac(current_stateSTATE_WR_CMD),
	.datad(WideOr13),
	.cin(gnd),
	.combout(src_startofpacket1),
	.cout());
defparam src_startofpacket.lut_mask = 16'hEAEE;
defparam src_startofpacket.sum_lutc_input = "datac";

cycloneive_lcell_comb \src_valid~0 (
	.dataa(stateST_IDLE),
	.datab(saved_grant_1),
	.datac(gnd),
	.datad(stateST_WAIT_RSP),
	.cin(gnd),
	.combout(src_valid),
	.cout());
defparam \src_valid~0 .lut_mask = 16'h0088;
defparam \src_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload[0]~1 (
	.dataa(stateST_SEND_HEADER),
	.datab(stateST_SEND_DATA_0),
	.datac(has_data_in),
	.datad(more_than_4bytes_data),
	.cin(gnd),
	.combout(src_payload_0),
	.cout());
defparam \src_payload[0]~1 .lut_mask = 16'h0ACE;
defparam \src_payload[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink0_ready~1 (
	.dataa(saved_grant_0),
	.datab(Selector18),
	.datac(stateST_SEND_DATA),
	.datad(\sink0_ready~0_combout ),
	.cin(gnd),
	.combout(sink0_ready),
	.cout());
defparam \sink0_ready~1 .lut_mask = 16'hA888;
defparam \sink0_ready~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[30]~3 (
	.dataa(saved_grant_1),
	.datab(csr_flash_cmd_wr_data_1_data_30),
	.datac(\src_data[30]~2_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(src_data_30),
	.cout());
defparam \src_data[30]~3 .lut_mask = 16'h88A0;
defparam \src_data[30]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[30]~5 (
	.dataa(mem_byteenable_reg_0),
	.datab(\src_data[30]~4_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_301),
	.cout());
defparam \src_data[30]~5 .lut_mask = 16'h8888;
defparam \src_data[30]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[30]~7 (
	.dataa(csr_control_data_7),
	.datab(current_stateSTATE_WR_DATA),
	.datac(\src_data[30]~6_combout ),
	.datad(cmd_valid1),
	.cin(gnd),
	.combout(src_data_302),
	.cout());
defparam \src_data[30]~7 .lut_mask = 16'hEAC0;
defparam \src_data[30]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[30]~8 (
	.dataa(src_data_30),
	.datab(saved_grant_0),
	.datac(src_data_302),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_303),
	.cout());
defparam \src_data[30]~8 .lut_mask = 16'hEAEA;
defparam \src_data[30]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[29]~10 (
	.dataa(saved_grant_1),
	.datab(csr_flash_cmd_wr_data_1_data_29),
	.datac(\src_data[29]~9_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(src_data_29),
	.cout());
defparam \src_data[29]~10 .lut_mask = 16'h88A0;
defparam \src_data[29]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[29]~12 (
	.dataa(csr_control_data_6),
	.datab(current_stateSTATE_WR_DATA),
	.datac(\src_data[29]~11_combout ),
	.datad(cmd_valid1),
	.cin(gnd),
	.combout(src_data_291),
	.cout());
defparam \src_data[29]~12 .lut_mask = 16'hEAC0;
defparam \src_data[29]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[29]~13 (
	.dataa(src_data_29),
	.datab(saved_grant_0),
	.datac(src_data_291),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_292),
	.cout());
defparam \src_data[29]~13 .lut_mask = 16'hEAEA;
defparam \src_data[29]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[28]~15 (
	.dataa(saved_grant_1),
	.datab(csr_flash_cmd_wr_data_1_data_28),
	.datac(\src_data[28]~14_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(src_data_28),
	.cout());
defparam \src_data[28]~15 .lut_mask = 16'h88A0;
defparam \src_data[28]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[28]~17 (
	.dataa(csr_control_data_5),
	.datab(current_stateSTATE_WR_DATA),
	.datac(\src_data[28]~16_combout ),
	.datad(cmd_valid1),
	.cin(gnd),
	.combout(src_data_281),
	.cout());
defparam \src_data[28]~17 .lut_mask = 16'hEAC0;
defparam \src_data[28]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[28]~18 (
	.dataa(src_data_28),
	.datab(saved_grant_0),
	.datac(src_data_281),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_282),
	.cout());
defparam \src_data[28]~18 .lut_mask = 16'hEAEA;
defparam \src_data[28]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[27]~20 (
	.dataa(saved_grant_1),
	.datab(csr_flash_cmd_wr_data_1_data_27),
	.datac(\src_data[27]~19_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(src_data_27),
	.cout());
defparam \src_data[27]~20 .lut_mask = 16'h88A0;
defparam \src_data[27]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[27]~22 (
	.dataa(csr_control_data_4),
	.datab(current_stateSTATE_WR_DATA),
	.datac(\src_data[27]~21_combout ),
	.datad(cmd_valid1),
	.cin(gnd),
	.combout(src_data_271),
	.cout());
defparam \src_data[27]~22 .lut_mask = 16'hEAC0;
defparam \src_data[27]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[27]~23 (
	.dataa(src_data_27),
	.datab(saved_grant_0),
	.datac(src_data_271),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_272),
	.cout());
defparam \src_data[27]~23 .lut_mask = 16'hEAEA;
defparam \src_data[27]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb WideOr1(
	.dataa(src_valid),
	.datab(saved_grant_0),
	.datac(cmd_valid),
	.datad(gnd),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hEAEA;
defparam WideOr1.sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload[0]~3 (
	.dataa(\src_payload[0]~2_combout ),
	.datab(saved_grant_1),
	.datac(stateST_SEND_DATA_1),
	.datad(src_payload_0),
	.cin(gnd),
	.combout(src_payload_01),
	.cout());
defparam \src_payload[0]~3 .lut_mask = 16'hEEEA;
defparam \src_payload[0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb sink1_ready(
	.dataa(saved_grant_1),
	.datab(Selector18),
	.datac(adap_out_cmd_ready),
	.datad(Selector181),
	.cin(gnd),
	.combout(sink1_ready1),
	.cout());
defparam sink1_ready.lut_mask = 16'hA888;
defparam sink1_ready.sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[11]~25 (
	.dataa(saved_grant_1),
	.datab(csr_flash_cmd_wr_data_1_data_11),
	.datac(\src_data[11]~24_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(src_data_11),
	.cout());
defparam \src_data[11]~25 .lut_mask = 16'h88A0;
defparam \src_data[11]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[11]~26 (
	.dataa(src_data_11),
	.datab(saved_grant_0),
	.datac(cmd_data_11),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_111),
	.cout());
defparam \src_data[11]~26 .lut_mask = 16'hEAEA;
defparam \src_data[11]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[18]~32 (
	.dataa(\src_data[18]~28_combout ),
	.datab(saved_grant_0),
	.datac(\src_data[18]~29_combout ),
	.datad(\src_data[18]~31_combout ),
	.cin(gnd),
	.combout(src_data_18),
	.cout());
defparam \src_data[18]~32 .lut_mask = 16'hEEEA;
defparam \src_data[18]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[19]~34 (
	.dataa(saved_grant_1),
	.datab(csr_flash_cmd_wr_data_1_data_19),
	.datac(\src_data[19]~33_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(src_data_19),
	.cout());
defparam \src_data[19]~34 .lut_mask = 16'h88A0;
defparam \src_data[19]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[19]~37 (
	.dataa(saved_grant_0),
	.datab(\src_data[19]~35_combout ),
	.datac(current_stateSTATE_WR_DATA),
	.datad(\src_data[19]~36_combout ),
	.cin(gnd),
	.combout(src_data_191),
	.cout());
defparam \src_data[19]~37 .lut_mask = 16'hA888;
defparam \src_data[19]~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[19]~38 (
	.dataa(src_data_19),
	.datab(src_data_191),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_192),
	.cout());
defparam \src_data[19]~38 .lut_mask = 16'hEEEE;
defparam \src_data[19]~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[21]~40 (
	.dataa(saved_grant_1),
	.datab(csr_flash_cmd_wr_data_1_data_21),
	.datac(\src_data[21]~39_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(src_data_21),
	.cout());
defparam \src_data[21]~40 .lut_mask = 16'h88A0;
defparam \src_data[21]~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[21]~43 (
	.dataa(is_burst_reg),
	.datab(mem_write_data_reg_21),
	.datac(\src_data[21]~41_combout ),
	.datad(\src_data[21]~42_combout ),
	.cin(gnd),
	.combout(src_data_211),
	.cout());
defparam \src_data[21]~43 .lut_mask = 16'hEAC0;
defparam \src_data[21]~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[21]~44 (
	.dataa(src_data_21),
	.datab(saved_grant_0),
	.datac(src_data_211),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_212),
	.cout());
defparam \src_data[21]~44 .lut_mask = 16'hEAEA;
defparam \src_data[21]~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[20]~46 (
	.dataa(saved_grant_1),
	.datab(csr_flash_cmd_wr_data_1_data_20),
	.datac(\src_data[20]~45_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(src_data_20),
	.cout());
defparam \src_data[20]~46 .lut_mask = 16'h88A0;
defparam \src_data[20]~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[20]~50 (
	.dataa(\src_data[20]~47_combout ),
	.datab(current_stateSTATE_WR_DATA),
	.datac(\src_data[20]~49_combout ),
	.datad(Selector20),
	.cin(gnd),
	.combout(src_data_201),
	.cout());
defparam \src_data[20]~50 .lut_mask = 16'h88B8;
defparam \src_data[20]~50 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[20]~51 (
	.dataa(src_data_20),
	.datab(saved_grant_0),
	.datac(src_data_201),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_202),
	.cout());
defparam \src_data[20]~51 .lut_mask = 16'hEAEA;
defparam \src_data[20]~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[22]~55 (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(\src_data[22]~53_combout ),
	.datad(\src_data[22]~54_combout ),
	.cin(gnd),
	.combout(src_data_22),
	.cout());
defparam \src_data[22]~55 .lut_mask = 16'hEAC0;
defparam \src_data[22]~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[23]~59 (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(\src_data[23]~57_combout ),
	.datad(\src_data[23]~58_combout ),
	.cin(gnd),
	.combout(src_data_23),
	.cout());
defparam \src_data[23]~59 .lut_mask = 16'hEAC0;
defparam \src_data[23]~59 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[24]~63 (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(\src_data[24]~61_combout ),
	.datad(\src_data[24]~62_combout ),
	.cin(gnd),
	.combout(src_data_24),
	.cout());
defparam \src_data[24]~63 .lut_mask = 16'hEAC0;
defparam \src_data[24]~63 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[25]~67 (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(\src_data[25]~65_combout ),
	.datad(\src_data[25]~66_combout ),
	.cin(gnd),
	.combout(src_data_25),
	.cout());
defparam \src_data[25]~67 .lut_mask = 16'hEAC0;
defparam \src_data[25]~67 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[26]~71 (
	.dataa(saved_grant_1),
	.datab(saved_grant_0),
	.datac(\src_data[26]~69_combout ),
	.datad(\src_data[26]~70_combout ),
	.cin(gnd),
	.combout(src_data_26),
	.cout());
defparam \src_data[26]~71 .lut_mask = 16'hEAC0;
defparam \src_data[26]~71 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[10]~73 (
	.dataa(saved_grant_1),
	.datab(\src_data[10]~72_combout ),
	.datac(csr_flash_cmd_wr_data_1_data_10),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(src_data_10),
	.cout());
defparam \src_data[10]~73 .lut_mask = 16'hA888;
defparam \src_data[10]~73 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[10]~74 (
	.dataa(src_data_10),
	.datab(saved_grant_0),
	.datac(cmd_data_10),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_101),
	.cout());
defparam \src_data[10]~74 .lut_mask = 16'hEAEA;
defparam \src_data[10]~74 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[8]~76 (
	.dataa(saved_grant_1),
	.datab(csr_flash_cmd_wr_data_1_data_8),
	.datac(\src_data[8]~75_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(src_data_8),
	.cout());
defparam \src_data[8]~76 .lut_mask = 16'h88A0;
defparam \src_data[8]~76 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[8]~77 (
	.dataa(src_data_8),
	.datab(saved_grant_0),
	.datac(cmd_data_8),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_81),
	.cout());
defparam \src_data[8]~77 .lut_mask = 16'hEAEA;
defparam \src_data[8]~77 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[13]~79 (
	.dataa(saved_grant_1),
	.datab(csr_flash_cmd_wr_data_1_data_13),
	.datac(\src_data[13]~78_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(src_data_13),
	.cout());
defparam \src_data[13]~79 .lut_mask = 16'h88A0;
defparam \src_data[13]~79 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[13]~80 (
	.dataa(src_data_13),
	.datab(saved_grant_0),
	.datac(cmd_data_13),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_131),
	.cout());
defparam \src_data[13]~80 .lut_mask = 16'hEAEA;
defparam \src_data[13]~80 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[17]~82 (
	.dataa(saved_grant_1),
	.datab(csr_flash_cmd_wr_data_1_data_17),
	.datac(\src_data[17]~81_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(src_data_17),
	.cout());
defparam \src_data[17]~82 .lut_mask = 16'h88A0;
defparam \src_data[17]~82 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[17]~84 (
	.dataa(\src_data[17]~83_combout ),
	.datab(csr_rd_inst_data_12),
	.datac(current_stateSTATE_READ_CMD),
	.datad(current_stateSTATE_WR_DATA),
	.cin(gnd),
	.combout(src_data_171),
	.cout());
defparam \src_data[17]~84 .lut_mask = 16'hAAC0;
defparam \src_data[17]~84 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[17]~85 (
	.dataa(src_data_17),
	.datab(saved_grant_0),
	.datac(src_data_171),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_172),
	.cout());
defparam \src_data[17]~85 .lut_mask = 16'hEAEA;
defparam \src_data[17]~85 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[16]~87 (
	.dataa(saved_grant_1),
	.datab(csr_flash_cmd_wr_data_1_data_16),
	.datac(\src_data[16]~86_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(src_data_16),
	.cout());
defparam \src_data[16]~87 .lut_mask = 16'h88A0;
defparam \src_data[16]~87 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[16]~89 (
	.dataa(\src_data[16]~88_combout ),
	.datab(csr_rd_inst_data_11),
	.datac(current_stateSTATE_READ_CMD),
	.datad(current_stateSTATE_WR_DATA),
	.cin(gnd),
	.combout(src_data_161),
	.cout());
defparam \src_data[16]~89 .lut_mask = 16'hAAC0;
defparam \src_data[16]~89 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[16]~90 (
	.dataa(src_data_16),
	.datab(saved_grant_0),
	.datac(src_data_161),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_162),
	.cout());
defparam \src_data[16]~90 .lut_mask = 16'hEAEA;
defparam \src_data[16]~90 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[15]~92 (
	.dataa(saved_grant_1),
	.datab(csr_flash_cmd_wr_data_1_data_15),
	.datac(\src_data[15]~91_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(src_data_15),
	.cout());
defparam \src_data[15]~92 .lut_mask = 16'h88A0;
defparam \src_data[15]~92 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[15]~93 (
	.dataa(src_data_15),
	.datab(saved_grant_0),
	.datac(cmd_data_15),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_151),
	.cout());
defparam \src_data[15]~93 .lut_mask = 16'hEAEA;
defparam \src_data[15]~93 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[14]~95 (
	.dataa(saved_grant_1),
	.datab(csr_flash_cmd_wr_data_1_data_14),
	.datac(\src_data[14]~94_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(src_data_14),
	.cout());
defparam \src_data[14]~95 .lut_mask = 16'h88A0;
defparam \src_data[14]~95 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[14]~96 (
	.dataa(src_data_14),
	.datab(saved_grant_0),
	.datac(cmd_data_14),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_141),
	.cout());
defparam \src_data[14]~96 .lut_mask = 16'hEAEA;
defparam \src_data[14]~96 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[9]~98 (
	.dataa(saved_grant_1),
	.datab(csr_flash_cmd_wr_data_1_data_9),
	.datac(\src_data[9]~97_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(src_data_9),
	.cout());
defparam \src_data[9]~98 .lut_mask = 16'h88A0;
defparam \src_data[9]~98 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[9]~99 (
	.dataa(src_data_9),
	.datab(saved_grant_0),
	.datac(cmd_data_9),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_91),
	.cout());
defparam \src_data[9]~99 .lut_mask = 16'hEAEA;
defparam \src_data[9]~99 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0]~102 (
	.dataa(\src_data[0]~101_combout ),
	.datab(\src_payload~4_combout ),
	.datac(\src_payload~5_combout ),
	.datad(cmd_data_0),
	.cin(gnd),
	.combout(src_data_0),
	.cout());
defparam \src_data[0]~102 .lut_mask = 16'hFEEE;
defparam \src_data[0]~102 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[4]~105 (
	.dataa(\src_data[4]~104_combout ),
	.datab(\src_payload~6_combout ),
	.datac(\src_payload~5_combout ),
	.datad(cmd_data_4),
	.cin(gnd),
	.combout(src_data_4),
	.cout());
defparam \src_data[4]~105 .lut_mask = 16'hFEEE;
defparam \src_data[4]~105 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[2]~108 (
	.dataa(\src_data[2]~107_combout ),
	.datab(\src_payload~7_combout ),
	.datac(cmd_data_2),
	.datad(\src_payload~5_combout ),
	.cin(gnd),
	.combout(src_data_2),
	.cout());
defparam \src_data[2]~108 .lut_mask = 16'hFEEE;
defparam \src_data[2]~108 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[1]~111 (
	.dataa(\src_data[1]~110_combout ),
	.datab(\src_payload~8_combout ),
	.datac(\src_payload~5_combout ),
	.datad(cmd_data_1),
	.cin(gnd),
	.combout(src_data_1),
	.cout());
defparam \src_data[1]~111 .lut_mask = 16'hFEEE;
defparam \src_data[1]~111 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[3]~114 (
	.dataa(\src_data[3]~113_combout ),
	.datab(\src_payload~9_combout ),
	.datac(\src_payload~5_combout ),
	.datad(cmd_data_3),
	.cin(gnd),
	.combout(src_data_3),
	.cout());
defparam \src_data[3]~114 .lut_mask = 16'hFEEE;
defparam \src_data[3]~114 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[5]~117 (
	.dataa(\src_data[5]~116_combout ),
	.datab(\src_payload~10_combout ),
	.datac(\src_payload~5_combout ),
	.datad(cmd_data_5),
	.cin(gnd),
	.combout(src_data_5),
	.cout());
defparam \src_data[5]~117 .lut_mask = 16'hFEEE;
defparam \src_data[5]~117 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[6]~120 (
	.dataa(\src_data[6]~119_combout ),
	.datab(\src_payload~11_combout ),
	.datac(\src_payload~5_combout ),
	.datad(cmd_data_6),
	.cin(gnd),
	.combout(src_data_6),
	.cout());
defparam \src_data[6]~120 .lut_mask = 16'hFEEE;
defparam \src_data[6]~120 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[7]~123 (
	.dataa(\src_data[7]~122_combout ),
	.datab(\src_payload~12_combout ),
	.datac(\src_payload~5_combout ),
	.datad(cmd_data_7),
	.cin(gnd),
	.combout(src_data_7),
	.cout());
defparam \src_data[7]~123 .lut_mask = 16'hFEEE;
defparam \src_data[7]~123 .sum_lutc_input = "datac";

cycloneive_lcell_comb \packet_in_progress~0 (
	.dataa(\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\packet_in_progress~0_combout ),
	.cout());
defparam \packet_in_progress~0 .lut_mask = 16'h5555;
defparam \packet_in_progress~0 .sum_lutc_input = "datac";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cycloneive_lcell_comb \update_grant~0 (
	.dataa(Selector182),
	.datab(src_payload_01),
	.datac(WideOr11),
	.datad(\packet_in_progress~q ),
	.cin(gnd),
	.combout(\update_grant~0_combout ),
	.cout());
defparam \update_grant~0 .lut_mask = 16'h808F;
defparam \update_grant~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~0 (
	.dataa(saved_grant_1),
	.datab(stateST_SEND_HEADER),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_payload~0_combout ),
	.cout());
defparam \src_payload~0 .lut_mask = 16'h8888;
defparam \src_payload~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink0_ready~0 (
	.dataa(Selector181),
	.datab(in_ready),
	.datac(WideOr01),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\sink0_ready~0_combout ),
	.cout());
defparam \sink0_ready~0 .lut_mask = 16'hAA80;
defparam \sink0_ready~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[30]~2 (
	.dataa(csr_flash_cmd_wr_data_0_data_30),
	.datab(csr_control_data_7),
	.datac(stateST_SEND_HEADER),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[30]~2_combout ),
	.cout());
defparam \src_data[30]~2 .lut_mask = 16'hAAC0;
defparam \src_data[30]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[30]~4 (
	.dataa(mem_byteenable_reg_3),
	.datab(mem_byteenable_reg_2),
	.datac(mem_byteenable_reg_1),
	.datad(is_burst_reg),
	.cin(gnd),
	.combout(\src_data[30]~4_combout ),
	.cout());
defparam \src_data[30]~4 .lut_mask = 16'h0080;
defparam \src_data[30]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[30]~6 (
	.dataa(is_burst_reg),
	.datab(mem_write_data_reg_30),
	.datac(src_data_301),
	.datad(out_payload_30),
	.cin(gnd),
	.combout(\src_data[30]~6_combout ),
	.cout());
defparam \src_data[30]~6 .lut_mask = 16'hEAC0;
defparam \src_data[30]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[29]~9 (
	.dataa(csr_flash_cmd_wr_data_0_data_29),
	.datab(csr_control_data_6),
	.datac(stateST_SEND_HEADER),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[29]~9_combout ),
	.cout());
defparam \src_data[29]~9 .lut_mask = 16'hAAC0;
defparam \src_data[29]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[29]~11 (
	.dataa(is_burst_reg),
	.datab(src_data_301),
	.datac(mem_write_data_reg_29),
	.datad(out_payload_29),
	.cin(gnd),
	.combout(\src_data[29]~11_combout ),
	.cout());
defparam \src_data[29]~11 .lut_mask = 16'hEAC0;
defparam \src_data[29]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[28]~14 (
	.dataa(csr_flash_cmd_wr_data_0_data_28),
	.datab(csr_control_data_5),
	.datac(stateST_SEND_HEADER),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[28]~14_combout ),
	.cout());
defparam \src_data[28]~14 .lut_mask = 16'hAAC0;
defparam \src_data[28]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[28]~16 (
	.dataa(is_burst_reg),
	.datab(src_data_301),
	.datac(mem_write_data_reg_28),
	.datad(out_payload_28),
	.cin(gnd),
	.combout(\src_data[28]~16_combout ),
	.cout());
defparam \src_data[28]~16 .lut_mask = 16'hEAC0;
defparam \src_data[28]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[27]~19 (
	.dataa(csr_flash_cmd_wr_data_0_data_27),
	.datab(csr_control_data_4),
	.datac(stateST_SEND_HEADER),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[27]~19_combout ),
	.cout());
defparam \src_data[27]~19 .lut_mask = 16'hAAC0;
defparam \src_data[27]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[27]~21 (
	.dataa(is_burst_reg),
	.datab(src_data_301),
	.datac(mem_write_data_reg_27),
	.datad(out_payload_27),
	.cin(gnd),
	.combout(\src_data[27]~21_combout ),
	.cout());
defparam \src_data[27]~21 .lut_mask = 16'hEAC0;
defparam \src_data[27]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload[0]~2 (
	.dataa(saved_grant_0),
	.datab(out_payload_32),
	.datac(current_stateSTATE_WR_DATA),
	.datad(WideOr13),
	.cin(gnd),
	.combout(\src_payload[0]~2_combout ),
	.cout());
defparam \src_payload[0]~2 .lut_mask = 16'h808A;
defparam \src_payload[0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[11]~24 (
	.dataa(csr_flash_cmd_wr_data_0_data_11),
	.datab(stateST_SEND_HEADER),
	.datac(has_data_out),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[11]~24_combout ),
	.cout());
defparam \src_data[11]~24 .lut_mask = 16'hAAC0;
defparam \src_data[11]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[18]~27 (
	.dataa(csr_flash_cmd_wr_data_0_data_18),
	.datab(stateST_SEND_HEADER),
	.datac(numb_data_0),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[18]~27_combout ),
	.cout());
defparam \src_data[18]~27 .lut_mask = 16'hAAC0;
defparam \src_data[18]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[18]~28 (
	.dataa(saved_grant_1),
	.datab(csr_flash_cmd_wr_data_1_data_18),
	.datac(\src_data[18]~27_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(\src_data[18]~28_combout ),
	.cout());
defparam \src_data[18]~28 .lut_mask = 16'h88A0;
defparam \src_data[18]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[18]~124 (
	.dataa(current_stateSTATE_WR_CMD),
	.datab(current_stateSTATE_READ_CMD),
	.datac(Add1),
	.datad(is_burst_reg),
	.cin(gnd),
	.combout(\src_data[18]~124_combout ),
	.cout());
defparam \src_data[18]~124 .lut_mask = 16'h00E0;
defparam \src_data[18]~124 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[18]~29 (
	.dataa(current_stateSTATE_STATUS_CMD),
	.datab(current_stateSTATE_POLL_CMD),
	.datac(\src_data[18]~124_combout ),
	.datad(current_stateSTATE_WR_DATA),
	.cin(gnd),
	.combout(\src_data[18]~29_combout ),
	.cout());
defparam \src_data[18]~29 .lut_mask = 16'h00FE;
defparam \src_data[18]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[18]~30 (
	.dataa(is_burst_reg),
	.datab(out_payload_18),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_data[18]~30_combout ),
	.cout());
defparam \src_data[18]~30 .lut_mask = 16'h8888;
defparam \src_data[18]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[18]~31 (
	.dataa(current_stateSTATE_WR_DATA),
	.datab(\src_data[18]~30_combout ),
	.datac(src_data_301),
	.datad(mem_write_data_reg_18),
	.cin(gnd),
	.combout(\src_data[18]~31_combout ),
	.cout());
defparam \src_data[18]~31 .lut_mask = 16'hA888;
defparam \src_data[18]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[19]~33 (
	.dataa(csr_flash_cmd_wr_data_0_data_19),
	.datab(stateST_SEND_HEADER),
	.datac(numb_data_1),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[19]~33_combout ),
	.cout());
defparam \src_data[19]~33 .lut_mask = 16'hAAC0;
defparam \src_data[19]~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[19]~35 (
	.dataa(Add11),
	.datab(current_stateSTATE_WR_DATA),
	.datac(is_burst_reg),
	.datad(Selector20),
	.cin(gnd),
	.combout(\src_data[19]~35_combout ),
	.cout());
defparam \src_data[19]~35 .lut_mask = 16'h0002;
defparam \src_data[19]~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[19]~36 (
	.dataa(is_burst_reg),
	.datab(src_data_301),
	.datac(mem_write_data_reg_19),
	.datad(out_payload_19),
	.cin(gnd),
	.combout(\src_data[19]~36_combout ),
	.cout());
defparam \src_data[19]~36 .lut_mask = 16'hEAC0;
defparam \src_data[19]~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[21]~39 (
	.dataa(csr_flash_cmd_wr_data_0_data_21),
	.datab(stateST_SEND_HEADER),
	.datac(numb_data_3),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[21]~39_combout ),
	.cout());
defparam \src_data[21]~39 .lut_mask = 16'hAAC0;
defparam \src_data[21]~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[21]~41 (
	.dataa(current_stateSTATE_WR_DATA),
	.datab(mem_byteenable_reg_0),
	.datac(\src_data[30]~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\src_data[21]~41_combout ),
	.cout());
defparam \src_data[21]~41 .lut_mask = 16'h8080;
defparam \src_data[21]~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[21]~42 (
	.dataa(out_payload_21),
	.datab(current_stateSTATE_WR_DATA),
	.datac(mem_burstcount_reg_1),
	.datad(Selector20),
	.cin(gnd),
	.combout(\src_data[21]~42_combout ),
	.cout());
defparam \src_data[21]~42 .lut_mask = 16'h88B8;
defparam \src_data[21]~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[20]~45 (
	.dataa(csr_flash_cmd_wr_data_0_data_20),
	.datab(stateST_SEND_HEADER),
	.datac(numb_data_2),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[20]~45_combout ),
	.cout());
defparam \src_data[20]~45 .lut_mask = 16'hAAC0;
defparam \src_data[20]~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[20]~47 (
	.dataa(is_burst_reg),
	.datab(src_data_301),
	.datac(mem_write_data_reg_20),
	.datad(out_payload_20),
	.cin(gnd),
	.combout(\src_data[20]~47_combout ),
	.cout());
defparam \src_data[20]~47 .lut_mask = 16'hEAC0;
defparam \src_data[20]~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[20]~48 (
	.dataa(mem_byteenable_reg_0),
	.datab(mem_byteenable_reg_3),
	.datac(mem_byteenable_reg_2),
	.datad(mem_byteenable_reg_1),
	.cin(gnd),
	.combout(\src_data[20]~48_combout ),
	.cout());
defparam \src_data[20]~48 .lut_mask = 16'h8000;
defparam \src_data[20]~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[20]~49 (
	.dataa(mem_burstcount_reg_0),
	.datab(\src_data[20]~48_combout ),
	.datac(gnd),
	.datad(is_burst_reg),
	.cin(gnd),
	.combout(\src_data[20]~49_combout ),
	.cout());
defparam \src_data[20]~49 .lut_mask = 16'hAACC;
defparam \src_data[20]~49 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[22]~52 (
	.dataa(out_payload_22),
	.datab(current_stateSTATE_WR_DATA),
	.datac(mem_burstcount_reg_2),
	.datad(Selector20),
	.cin(gnd),
	.combout(\src_data[22]~52_combout ),
	.cout());
defparam \src_data[22]~52 .lut_mask = 16'h88B8;
defparam \src_data[22]~52 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[22]~53 (
	.dataa(is_burst_reg),
	.datab(\src_data[21]~41_combout ),
	.datac(mem_write_data_reg_22),
	.datad(\src_data[22]~52_combout ),
	.cin(gnd),
	.combout(\src_data[22]~53_combout ),
	.cout());
defparam \src_data[22]~53 .lut_mask = 16'hEAC0;
defparam \src_data[22]~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[22]~54 (
	.dataa(csr_flash_cmd_wr_data_0_data_22),
	.datab(csr_flash_cmd_wr_data_1_data_22),
	.datac(stateST_SEND_DATA_1),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[22]~54_combout ),
	.cout());
defparam \src_data[22]~54 .lut_mask = 16'hEAC0;
defparam \src_data[22]~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[23]~56 (
	.dataa(out_payload_23),
	.datab(current_stateSTATE_WR_DATA),
	.datac(mem_burstcount_reg_3),
	.datad(Selector20),
	.cin(gnd),
	.combout(\src_data[23]~56_combout ),
	.cout());
defparam \src_data[23]~56 .lut_mask = 16'h88B8;
defparam \src_data[23]~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[23]~57 (
	.dataa(is_burst_reg),
	.datab(\src_data[21]~41_combout ),
	.datac(mem_write_data_reg_23),
	.datad(\src_data[23]~56_combout ),
	.cin(gnd),
	.combout(\src_data[23]~57_combout ),
	.cout());
defparam \src_data[23]~57 .lut_mask = 16'hEAC0;
defparam \src_data[23]~57 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[23]~58 (
	.dataa(csr_flash_cmd_wr_data_0_data_23),
	.datab(csr_flash_cmd_wr_data_1_data_23),
	.datac(stateST_SEND_DATA_1),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[23]~58_combout ),
	.cout());
defparam \src_data[23]~58 .lut_mask = 16'hEAC0;
defparam \src_data[23]~58 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[24]~60 (
	.dataa(out_payload_24),
	.datab(current_stateSTATE_WR_DATA),
	.datac(mem_burstcount_reg_4),
	.datad(Selector20),
	.cin(gnd),
	.combout(\src_data[24]~60_combout ),
	.cout());
defparam \src_data[24]~60 .lut_mask = 16'h88B8;
defparam \src_data[24]~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[24]~61 (
	.dataa(is_burst_reg),
	.datab(\src_data[21]~41_combout ),
	.datac(mem_write_data_reg_24),
	.datad(\src_data[24]~60_combout ),
	.cin(gnd),
	.combout(\src_data[24]~61_combout ),
	.cout());
defparam \src_data[24]~61 .lut_mask = 16'hEAC0;
defparam \src_data[24]~61 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[24]~62 (
	.dataa(csr_flash_cmd_wr_data_0_data_24),
	.datab(csr_flash_cmd_wr_data_1_data_24),
	.datac(stateST_SEND_DATA_1),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[24]~62_combout ),
	.cout());
defparam \src_data[24]~62 .lut_mask = 16'hEAC0;
defparam \src_data[24]~62 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[25]~64 (
	.dataa(out_payload_25),
	.datab(current_stateSTATE_WR_DATA),
	.datac(mem_burstcount_reg_5),
	.datad(Selector20),
	.cin(gnd),
	.combout(\src_data[25]~64_combout ),
	.cout());
defparam \src_data[25]~64 .lut_mask = 16'h88B8;
defparam \src_data[25]~64 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[25]~65 (
	.dataa(is_burst_reg),
	.datab(\src_data[21]~41_combout ),
	.datac(mem_write_data_reg_25),
	.datad(\src_data[25]~64_combout ),
	.cin(gnd),
	.combout(\src_data[25]~65_combout ),
	.cout());
defparam \src_data[25]~65 .lut_mask = 16'hEAC0;
defparam \src_data[25]~65 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[25]~66 (
	.dataa(csr_flash_cmd_wr_data_0_data_25),
	.datab(csr_flash_cmd_wr_data_1_data_25),
	.datac(stateST_SEND_DATA_1),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[25]~66_combout ),
	.cout());
defparam \src_data[25]~66 .lut_mask = 16'hEAC0;
defparam \src_data[25]~66 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[26]~68 (
	.dataa(out_payload_26),
	.datab(current_stateSTATE_WR_DATA),
	.datac(mem_burstcount_reg_6),
	.datad(Selector20),
	.cin(gnd),
	.combout(\src_data[26]~68_combout ),
	.cout());
defparam \src_data[26]~68 .lut_mask = 16'h88B8;
defparam \src_data[26]~68 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[26]~69 (
	.dataa(is_burst_reg),
	.datab(\src_data[21]~41_combout ),
	.datac(mem_write_data_reg_26),
	.datad(\src_data[26]~68_combout ),
	.cin(gnd),
	.combout(\src_data[26]~69_combout ),
	.cout());
defparam \src_data[26]~69 .lut_mask = 16'hEAC0;
defparam \src_data[26]~69 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[26]~70 (
	.dataa(csr_flash_cmd_wr_data_0_data_26),
	.datab(csr_flash_cmd_wr_data_1_data_26),
	.datac(stateST_SEND_DATA_1),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[26]~70_combout ),
	.cout());
defparam \src_data[26]~70 .lut_mask = 16'hEAC0;
defparam \src_data[26]~70 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[10]~72 (
	.dataa(csr_flash_cmd_wr_data_0_data_10),
	.datab(Selector34),
	.datac(stateST_SEND_DATA_0),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(\src_data[10]~72_combout ),
	.cout());
defparam \src_data[10]~72 .lut_mask = 16'h00AC;
defparam \src_data[10]~72 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[8]~75 (
	.dataa(csr_flash_cmd_wr_data_0_data_8),
	.datab(stateST_SEND_HEADER),
	.datac(has_addr),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[8]~75_combout ),
	.cout());
defparam \src_data[8]~75 .lut_mask = 16'hAAC0;
defparam \src_data[8]~75 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[13]~78 (
	.dataa(csr_flash_cmd_wr_data_0_data_13),
	.datab(stateST_SEND_HEADER),
	.datac(numb_dummy_0),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[13]~78_combout ),
	.cout());
defparam \src_data[13]~78 .lut_mask = 16'hAAC0;
defparam \src_data[13]~78 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[17]~81 (
	.dataa(csr_flash_cmd_wr_data_0_data_17),
	.datab(stateST_SEND_HEADER),
	.datac(numb_dummy_4),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[17]~81_combout ),
	.cout());
defparam \src_data[17]~81 .lut_mask = 16'hAAC0;
defparam \src_data[17]~81 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[17]~83 (
	.dataa(is_burst_reg),
	.datab(src_data_301),
	.datac(mem_write_data_reg_17),
	.datad(out_payload_17),
	.cin(gnd),
	.combout(\src_data[17]~83_combout ),
	.cout());
defparam \src_data[17]~83 .lut_mask = 16'hEAC0;
defparam \src_data[17]~83 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[16]~86 (
	.dataa(csr_flash_cmd_wr_data_0_data_16),
	.datab(stateST_SEND_HEADER),
	.datac(numb_dummy_3),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[16]~86_combout ),
	.cout());
defparam \src_data[16]~86 .lut_mask = 16'hAAC0;
defparam \src_data[16]~86 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[16]~88 (
	.dataa(is_burst_reg),
	.datab(src_data_301),
	.datac(mem_write_data_reg_16),
	.datad(out_payload_16),
	.cin(gnd),
	.combout(\src_data[16]~88_combout ),
	.cout());
defparam \src_data[16]~88 .lut_mask = 16'hEAC0;
defparam \src_data[16]~88 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[15]~91 (
	.dataa(csr_flash_cmd_wr_data_0_data_15),
	.datab(stateST_SEND_HEADER),
	.datac(numb_dummy_2),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[15]~91_combout ),
	.cout());
defparam \src_data[15]~91 .lut_mask = 16'hAAC0;
defparam \src_data[15]~91 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[14]~94 (
	.dataa(csr_flash_cmd_wr_data_0_data_14),
	.datab(stateST_SEND_HEADER),
	.datac(numb_dummy_1),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[14]~94_combout ),
	.cout());
defparam \src_data[14]~94 .lut_mask = 16'hAAC0;
defparam \src_data[14]~94 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[9]~97 (
	.dataa(csr_flash_cmd_wr_data_0_data_9),
	.datab(stateST_SEND_HEADER),
	.datac(is_4bytes_addr),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[9]~97_combout ),
	.cout());
defparam \src_data[9]~97 .lut_mask = 16'hAAC0;
defparam \src_data[9]~97 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0]~100 (
	.dataa(csr_flash_cmd_wr_data_0_data_0),
	.datab(stateST_SEND_HEADER),
	.datac(opcode_0),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[0]~100_combout ),
	.cout());
defparam \src_data[0]~100 .lut_mask = 16'hAAC0;
defparam \src_data[0]~100 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0]~101 (
	.dataa(saved_grant_1),
	.datab(csr_flash_cmd_wr_data_1_data_0),
	.datac(\src_data[0]~100_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(\src_data[0]~101_combout ),
	.cout());
defparam \src_data[0]~101 .lut_mask = 16'h88A0;
defparam \src_data[0]~101 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~4 (
	.dataa(saved_grant_0),
	.datab(current_stateSTATE_WR_DATA),
	.datac(is_burst_reg),
	.datad(out_payload_0),
	.cin(gnd),
	.combout(\src_payload~4_combout ),
	.cout());
defparam \src_payload~4 .lut_mask = 16'h8000;
defparam \src_payload~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~5 (
	.dataa(saved_grant_0),
	.datab(gnd),
	.datac(current_stateSTATE_WR_DATA),
	.datad(is_burst_reg),
	.cin(gnd),
	.combout(\src_payload~5_combout ),
	.cout());
defparam \src_payload~5 .lut_mask = 16'h0AAA;
defparam \src_payload~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[4]~103 (
	.dataa(csr_flash_cmd_wr_data_0_data_4),
	.datab(stateST_SEND_HEADER),
	.datac(opcode_4),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[4]~103_combout ),
	.cout());
defparam \src_data[4]~103 .lut_mask = 16'hAAC0;
defparam \src_data[4]~103 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[4]~104 (
	.dataa(saved_grant_1),
	.datab(csr_flash_cmd_wr_data_1_data_4),
	.datac(\src_data[4]~103_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(\src_data[4]~104_combout ),
	.cout());
defparam \src_data[4]~104 .lut_mask = 16'h88A0;
defparam \src_data[4]~104 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~6 (
	.dataa(saved_grant_0),
	.datab(current_stateSTATE_WR_DATA),
	.datac(is_burst_reg),
	.datad(out_payload_4),
	.cin(gnd),
	.combout(\src_payload~6_combout ),
	.cout());
defparam \src_payload~6 .lut_mask = 16'h8000;
defparam \src_payload~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[2]~106 (
	.dataa(csr_flash_cmd_wr_data_0_data_2),
	.datab(stateST_SEND_HEADER),
	.datac(opcode_2),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[2]~106_combout ),
	.cout());
defparam \src_data[2]~106 .lut_mask = 16'hAAC0;
defparam \src_data[2]~106 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[2]~107 (
	.dataa(saved_grant_1),
	.datab(csr_flash_cmd_wr_data_1_data_2),
	.datac(\src_data[2]~106_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(\src_data[2]~107_combout ),
	.cout());
defparam \src_data[2]~107 .lut_mask = 16'h88A0;
defparam \src_data[2]~107 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~7 (
	.dataa(saved_grant_0),
	.datab(current_stateSTATE_WR_DATA),
	.datac(is_burst_reg),
	.datad(out_payload_2),
	.cin(gnd),
	.combout(\src_payload~7_combout ),
	.cout());
defparam \src_payload~7 .lut_mask = 16'h8000;
defparam \src_payload~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[1]~109 (
	.dataa(csr_flash_cmd_wr_data_0_data_1),
	.datab(stateST_SEND_HEADER),
	.datac(opcode_1),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[1]~109_combout ),
	.cout());
defparam \src_data[1]~109 .lut_mask = 16'hAAC0;
defparam \src_data[1]~109 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[1]~110 (
	.dataa(saved_grant_1),
	.datab(csr_flash_cmd_wr_data_1_data_1),
	.datac(\src_data[1]~109_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(\src_data[1]~110_combout ),
	.cout());
defparam \src_data[1]~110 .lut_mask = 16'h88A0;
defparam \src_data[1]~110 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~8 (
	.dataa(saved_grant_0),
	.datab(current_stateSTATE_WR_DATA),
	.datac(is_burst_reg),
	.datad(out_payload_1),
	.cin(gnd),
	.combout(\src_payload~8_combout ),
	.cout());
defparam \src_payload~8 .lut_mask = 16'h8000;
defparam \src_payload~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[3]~112 (
	.dataa(csr_flash_cmd_wr_data_0_data_3),
	.datab(stateST_SEND_HEADER),
	.datac(opcode_3),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[3]~112_combout ),
	.cout());
defparam \src_data[3]~112 .lut_mask = 16'hAAC0;
defparam \src_data[3]~112 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[3]~113 (
	.dataa(saved_grant_1),
	.datab(csr_flash_cmd_wr_data_1_data_3),
	.datac(\src_data[3]~112_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(\src_data[3]~113_combout ),
	.cout());
defparam \src_data[3]~113 .lut_mask = 16'h88A0;
defparam \src_data[3]~113 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~9 (
	.dataa(saved_grant_0),
	.datab(current_stateSTATE_WR_DATA),
	.datac(is_burst_reg),
	.datad(out_payload_3),
	.cin(gnd),
	.combout(\src_payload~9_combout ),
	.cout());
defparam \src_payload~9 .lut_mask = 16'h8000;
defparam \src_payload~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[5]~115 (
	.dataa(csr_flash_cmd_wr_data_0_data_5),
	.datab(stateST_SEND_HEADER),
	.datac(opcode_5),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[5]~115_combout ),
	.cout());
defparam \src_data[5]~115 .lut_mask = 16'hAAC0;
defparam \src_data[5]~115 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[5]~116 (
	.dataa(saved_grant_1),
	.datab(csr_flash_cmd_wr_data_1_data_5),
	.datac(\src_data[5]~115_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(\src_data[5]~116_combout ),
	.cout());
defparam \src_data[5]~116 .lut_mask = 16'h88A0;
defparam \src_data[5]~116 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~10 (
	.dataa(saved_grant_0),
	.datab(current_stateSTATE_WR_DATA),
	.datac(is_burst_reg),
	.datad(out_payload_5),
	.cin(gnd),
	.combout(\src_payload~10_combout ),
	.cout());
defparam \src_payload~10 .lut_mask = 16'h8000;
defparam \src_payload~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[6]~118 (
	.dataa(csr_flash_cmd_wr_data_0_data_6),
	.datab(stateST_SEND_HEADER),
	.datac(opcode_6),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[6]~118_combout ),
	.cout());
defparam \src_data[6]~118 .lut_mask = 16'hAAC0;
defparam \src_data[6]~118 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[6]~119 (
	.dataa(saved_grant_1),
	.datab(csr_flash_cmd_wr_data_1_data_6),
	.datac(\src_data[6]~118_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(\src_data[6]~119_combout ),
	.cout());
defparam \src_data[6]~119 .lut_mask = 16'h88A0;
defparam \src_data[6]~119 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~11 (
	.dataa(saved_grant_0),
	.datab(current_stateSTATE_WR_DATA),
	.datac(is_burst_reg),
	.datad(out_payload_6),
	.cin(gnd),
	.combout(\src_payload~11_combout ),
	.cout());
defparam \src_payload~11 .lut_mask = 16'h8000;
defparam \src_payload~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[7]~121 (
	.dataa(csr_flash_cmd_wr_data_0_data_7),
	.datab(stateST_SEND_HEADER),
	.datac(opcode_7),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\src_data[7]~121_combout ),
	.cout());
defparam \src_data[7]~121 .lut_mask = 16'hAAC0;
defparam \src_data[7]~121 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[7]~122 (
	.dataa(saved_grant_1),
	.datab(csr_flash_cmd_wr_data_1_data_7),
	.datac(\src_data[7]~121_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(\src_data[7]~122_combout ),
	.cout());
defparam \src_data[7]~122 .lut_mask = 16'h88A0;
defparam \src_data[7]~122 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload~12 (
	.dataa(saved_grant_0),
	.datab(current_stateSTATE_WR_DATA),
	.datac(is_burst_reg),
	.datad(out_payload_7),
	.cin(gnd),
	.combout(\src_payload~12_combout ),
	.cout());
defparam \src_payload~12 .lut_mask = 16'h8000;
defparam \src_payload~12 .sum_lutc_input = "datac";

endmodule

module flashLoader_altera_merlin_arbitrator (
	stateST_IDLE,
	stateST_WAIT_RSP,
	cmd_valid,
	grant_1)/* synthesis synthesis_greybox=0 */;
input 	stateST_IDLE;
input 	stateST_WAIT_RSP;
input 	cmd_valid;
output 	grant_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \grant[1]~0 (
	.dataa(stateST_WAIT_RSP),
	.datab(cmd_valid),
	.datac(gnd),
	.datad(stateST_IDLE),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~0 .lut_mask = 16'h1100;
defparam \grant[1]~0 .sum_lutc_input = "datac";

endmodule

module flashLoader_flashLoader_intel_generic_serial_flash_interface_top_0_qspi_inf_inst (
	data_num_lines_1,
	data_num_lines_2,
	addr_num_lines_2,
	addr_num_lines_1,
	flash_clk_reg1,
	oe_reg1,
	ncs_reg_0,
	flash_data_out_reg_0,
	csr_delay_setting_data_0,
	csr_clk_baud_rate_data_0,
	qspi_interface_en,
	csr_rd_capturing_data_0,
	altera_reset_synchronizer_int_chain_out,
	csr_delay_setting_data_1,
	csr_clk_baud_rate_data_1,
	csr_rd_capturing_data_1,
	csr_delay_setting_data_2,
	csr_clk_baud_rate_data_2,
	csr_rd_capturing_data_2,
	csr_delay_setting_data_3,
	csr_clk_baud_rate_data_3,
	csr_rd_capturing_data_3,
	csr_delay_setting_data_4,
	csr_clk_baud_rate_data_4,
	csr_delay_setting_data_5,
	csr_delay_setting_data_6,
	csr_delay_setting_data_7,
	in_cmd_channel_reg_1,
	in_cmd_channel_reg_0,
	header_information_30,
	header_information_29,
	header_information_28,
	header_information_27,
	stateST_IDLE,
	stateST_SEND_DATA,
	stateST_SEND_ADDR,
	op_num_lines_1,
	data_num_lines_0,
	op_num_lines_0,
	WideOr0,
	in_ready,
	op_num_lines_2,
	WideOr01,
	header_information_11,
	stateST_SEND_OPCODE,
	Selector8,
	demux_channel_2,
	in_cmd_ready,
	addr_num_lines_0,
	WideOr02,
	out_rsp_valid1,
	WideOr03,
	WideOr04,
	WideOr05,
	out_rsp_data_0,
	out_rsp_data_1,
	out_rsp_data_2,
	out_rsp_data_3,
	out_rsp_data_4,
	out_rsp_data_5,
	out_rsp_data_6,
	out_rsp_data_7,
	header_information_13,
	header_information_17,
	header_information_16,
	header_information_15,
	header_information_14,
	WideOr06,
	Selector20,
	Selector16,
	Selector12,
	Selector14,
	Selector15,
	Selector13,
	Selector11,
	Selector10,
	Selector9,
	Selector17,
	clk_clk,
	dut_asmiblock)/* synthesis synthesis_greybox=0 */;
input 	data_num_lines_1;
input 	data_num_lines_2;
input 	addr_num_lines_2;
input 	addr_num_lines_1;
output 	flash_clk_reg1;
output 	oe_reg1;
output 	ncs_reg_0;
output 	flash_data_out_reg_0;
input 	csr_delay_setting_data_0;
input 	csr_clk_baud_rate_data_0;
input 	qspi_interface_en;
input 	csr_rd_capturing_data_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	csr_delay_setting_data_1;
input 	csr_clk_baud_rate_data_1;
input 	csr_rd_capturing_data_1;
input 	csr_delay_setting_data_2;
input 	csr_clk_baud_rate_data_2;
input 	csr_rd_capturing_data_2;
input 	csr_delay_setting_data_3;
input 	csr_clk_baud_rate_data_3;
input 	csr_rd_capturing_data_3;
input 	csr_delay_setting_data_4;
input 	csr_clk_baud_rate_data_4;
input 	csr_delay_setting_data_5;
input 	csr_delay_setting_data_6;
input 	csr_delay_setting_data_7;
input 	in_cmd_channel_reg_1;
input 	in_cmd_channel_reg_0;
input 	header_information_30;
input 	header_information_29;
input 	header_information_28;
input 	header_information_27;
input 	stateST_IDLE;
input 	stateST_SEND_DATA;
input 	stateST_SEND_ADDR;
input 	op_num_lines_1;
input 	data_num_lines_0;
input 	op_num_lines_0;
output 	WideOr0;
output 	in_ready;
input 	op_num_lines_2;
output 	WideOr01;
input 	header_information_11;
input 	stateST_SEND_OPCODE;
input 	Selector8;
output 	demux_channel_2;
output 	in_cmd_ready;
input 	addr_num_lines_0;
output 	WideOr02;
output 	out_rsp_valid1;
output 	WideOr03;
output 	WideOr04;
output 	WideOr05;
output 	out_rsp_data_0;
output 	out_rsp_data_1;
output 	out_rsp_data_2;
output 	out_rsp_data_3;
output 	out_rsp_data_4;
output 	out_rsp_data_5;
output 	out_rsp_data_6;
output 	out_rsp_data_7;
input 	header_information_13;
input 	header_information_17;
input 	header_information_16;
input 	header_information_15;
input 	header_information_14;
output 	WideOr06;
input 	Selector20;
input 	Selector16;
input 	Selector12;
input 	Selector14;
input 	Selector15;
input 	Selector13;
input 	Selector11;
input 	Selector10;
input 	Selector9;
input 	Selector17;
input 	clk_clk;
input 	dut_asmiblock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \WideOr7~0_combout ;
wire \clk_div_new_inst_2|clk_track~q ;
wire \clk_div_new_inst_2|clk_out~0_combout ;
wire \inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|out_payload[12]~q ;
wire \inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|out_payload[2]~q ;
wire \inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|out_payload[1]~q ;
wire \inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|out_payload[0]~q ;
wire \adapter_8_4_inst|out_valid~q ;
wire \qspi_inf_mux_inst|qspi_inf_mux|arb|grant[0]~2_combout ;
wire \adapter_8_1_inst|out_valid~q ;
wire \adapter_8_2_inst|out_valid~q ;
wire \qspi_inf_mux_inst|qspi_inf_mux|request[1]~combout ;
wire \qspi_inf_mux_inst|qspi_inf_mux|arb|adder|full_adder.cout[1]~combout ;
wire \qspi_inf_mux_inst|qspi_inf_mux|arb|adder|cout~0_combout ;
wire \inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|mem_used[9]~q ;
wire \adapter_8_1_inst|in_ready~combout ;
wire \adapter_8_2_inst|state_register[1]~q ;
wire \adapter_8_2_inst|state_register[0]~q ;
wire \adapter_8_2_inst|a_valid~q ;
wire \qspi_inf_mux_inst|qspi_inf_mux|arb|adder|sum[1]~combout ;
wire \qspi_inf_mux_inst|qspi_inf_mux|request[2]~combout ;
wire \qspi_inf_mux_inst|qspi_inf_mux|arb|adder|cout~1_combout ;
wire \adapter_8_2_inst|always4~1_combout ;
wire \adapter_8_4_inst|state_register[0]~q ;
wire \adapter_8_4_inst|always4~0_combout ;
wire \adapter_8_4_inst|always4~1_combout ;
wire \adapter_8_4_inst|a_valid~q ;
wire \inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|out_valid~q ;
wire \clk_div_new_inst_2|Equal0~1_combout ;
wire \clk_div_new_inst_2|Equal0~2_combout ;
wire \clk_div_new_inst_2|enable_d~q ;
wire \clk_div_new_inst_2|Add1~1_combout ;
wire \inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|out_payload[16]~q ;
wire \inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|out_payload[8]~q ;
wire \WideOr7~combout ;
wire \clk_div_new_inst_2|Equal0~3_combout ;
wire \adapter_8_2_inst|in_ready~combout ;
wire \demux_channel[1]~2_combout ;
wire \demux_channel[1]~3_combout ;
wire \demux_channel[0]~4_combout ;
wire \demux_channel[0]~5_combout ;
wire \qspi_inf_mux_inst|qspi_inf_mux|arb|grant[0]~3_combout ;
wire \qspi_inf_mux_inst|qspi_inf_mux|WideOr1~2_combout ;
wire \inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|write~0_combout ;
wire \adapter_8_4_inst|out_endofpacket~q ;
wire \adapter_8_1_inst|out_endofpacket~q ;
wire \adapter_8_2_inst|out_endofpacket~q ;
wire \qspi_inf_mux_inst|qspi_inf_mux|src_payload[0]~1_combout ;
wire \demux_channel[2]~6_combout ;
wire \demultiplexer_inst|src0_valid~combout ;
wire \demultiplexer_inst|src1_valid~combout ;
wire \demultiplexer_inst|src2_valid~combout ;
wire \adapter_8_4_inst|out_data[0]~q ;
wire \adapter_8_1_inst|out_data[0]~q ;
wire \adapter_8_2_inst|out_data[0]~q ;
wire \qspi_inf_mux_inst|qspi_inf_mux|src_data[0]~1_combout ;
wire \adapter_8_4_inst|out_channel[2]~q ;
wire \adapter_8_1_inst|out_channel[2]~q ;
wire \adapter_8_2_inst|out_channel[2]~q ;
wire \qspi_inf_mux_inst|qspi_inf_mux|src_channel[2]~1_combout ;
wire \adapter_8_4_inst|out_channel[1]~q ;
wire \adapter_8_1_inst|out_channel[1]~q ;
wire \adapter_8_2_inst|out_channel[1]~q ;
wire \qspi_inf_mux_inst|qspi_inf_mux|src_channel[1]~3_combout ;
wire \adapter_8_4_inst|out_channel[0]~q ;
wire \adapter_8_1_inst|out_channel[0]~q ;
wire \adapter_8_2_inst|out_channel[0]~q ;
wire \qspi_inf_mux_inst|qspi_inf_mux|src_channel[0]~5_combout ;
wire \adapter_8_4_inst|out_channel[8]~q ;
wire \adapter_8_1_inst|out_channel[8]~q ;
wire \adapter_8_2_inst|out_channel[8]~q ;
wire \qspi_inf_mux_inst|qspi_inf_mux|src_channel[8]~7_combout ;
wire \clk_div_new_inst_2|rising_edge~combout ;
wire \Selector0~0_combout ;
wire \state.ST_IDLE~q ;
wire \LessThan0~0_combout ;
wire \Equal14~1_combout ;
wire \cs_assert_cnt_next~4_combout ;
wire \cs_assert_cnt[1]~q ;
wire \Equal14~2_combout ;
wire \cs_assert_cnt_next~3_combout ;
wire \cs_assert_cnt[0]~q ;
wire \cs_assert_cnt_next~5_combout ;
wire \cs_assert_cnt[2]~q ;
wire \Add3~0_combout ;
wire \cs_assert_cnt_next~2_combout ;
wire \cs_assert_cnt[3]~q ;
wire \Equal14~0_combout ;
wire \Equal14~3_combout ;
wire \ncs_wire[0]~2_combout ;
wire \Selector1~0_combout ;
wire \state.ST_ASSERT_CS_DLY~q ;
wire \Selector2~0_combout ;
wire \state.ST_START_CLK~q ;
wire \require_rdata_reg~0_combout ;
wire \require_rdata_reg~q ;
wire \state.ST_ASSERT_CS~q ;
wire \fifo_pop_out~0_combout ;
wire \fifo_pop_out~1_combout ;
wire \next_state~1_combout ;
wire \Selector3~0_combout ;
wire \state.ST_SEND~q ;
wire \next_state~0_combout ;
wire \LessThan1~0_combout ;
wire \Selector5~0_combout ;
wire \Selector5~1_combout ;
wire \next_state~2_combout ;
wire \Add0~1 ;
wire \Add0~3 ;
wire \Add0~5 ;
wire \Add0~7 ;
wire \Add0~8_combout ;
wire \dummy_cnt[0]~5_combout ;
wire \always6~1_combout ;
wire \dummy_cnt[0]~q ;
wire \dummy_cnt[0]~6 ;
wire \dummy_cnt[1]~7_combout ;
wire \dummy_cnt[1]~q ;
wire \dummy_cnt[1]~8 ;
wire \dummy_cnt[2]~9_combout ;
wire \dummy_cnt[2]~q ;
wire \dummy_cnt[2]~10 ;
wire \dummy_cnt[3]~11_combout ;
wire \dummy_cnt[3]~q ;
wire \dummy_cnt[3]~12 ;
wire \dummy_cnt[4]~13_combout ;
wire \dummy_cnt[4]~q ;
wire \Add0~4_combout ;
wire \Add0~6_combout ;
wire \dummy_cnt_done~0_combout ;
wire \Add0~0_combout ;
wire \Add0~2_combout ;
wire \dummy_cnt_done~1_combout ;
wire \dummy_cnt_done~2_combout ;
wire \dummy_cnt_done~3_combout ;
wire \Selector4~0_combout ;
wire \state.ST_DUMMY_CYCLES~q ;
wire \Selector5~2_combout ;
wire \state.ST_RECEIVE~q ;
wire \Selector6~0_combout ;
wire \Selector6~1_combout ;
wire \state.ST_STOP_CLK~q ;
wire \cs_deassert_cnt_next~4_combout ;
wire \cs_deassert_cnt[1]~q ;
wire \Add5~0_combout ;
wire \cs_deassert_cnt_next~5_combout ;
wire \cs_deassert_cnt[3]~q ;
wire \Equal15~1_combout ;
wire \Equal15~2_combout ;
wire \cs_deassert_cnt_next~7_combout ;
wire \cs_deassert_cnt[0]~q ;
wire \cs_deassert_cnt_next~6_combout ;
wire \cs_deassert_cnt[2]~q ;
wire \Equal15~0_combout ;
wire \Equal15~3_combout ;
wire \Selector7~0_combout ;
wire \Selector8~0_combout ;
wire \state.ST_DEASSERT_CS_DLY~q ;
wire \Selector7~1_combout ;
wire \state.ST_DEASSERT_CS~q ;
wire \ncs_wire[0]~0_combout ;
wire \ncs_wire[0]~1_combout ;
wire \ncs_wire[0]~3_combout ;
wire \flash_data_out[0]~0_combout ;
wire \demux_channel[2]~0_combout ;
wire \Equal0~0_combout ;
wire \read_capture_delay_reg[0]~q ;
wire \read_capture_delay_reg~9_combout ;
wire \read_capture_delay_reg[1]~q ;
wire \read_capture_delay_reg~8_combout ;
wire \read_capture_delay_reg[2]~q ;
wire \read_capture_delay_reg~10_combout ;
wire \read_capture_delay_reg[3]~q ;
wire \read_capture_delay_reg~6_combout ;
wire \read_capture_delay_reg[4]~q ;
wire \read_capture_delay_reg~4_combout ;
wire \read_capture_delay_reg[5]~q ;
wire \read_capture_delay_reg~5_combout ;
wire \read_capture_delay_reg[6]~q ;
wire \read_capture_delay_reg~7_combout ;
wire \read_capture_delay_reg[7]~q ;
wire \read_capture_delay_reg~2_combout ;
wire \read_capture_delay_reg[8]~q ;
wire \read_capture_delay_reg~1_combout ;
wire \read_capture_delay_reg[9]~q ;
wire \read_capture_delay_reg~0_combout ;
wire \read_capture_delay_reg[10]~q ;
wire \Mux0~0_combout ;
wire \read_capture_delay_reg~3_combout ;
wire \read_capture_delay_reg[11]~q ;
wire \Mux0~1_combout ;
wire \Mux0~2_combout ;
wire \Mux0~3_combout ;
wire \Mux0~4_combout ;
wire \Mux0~5_combout ;
wire \Mux0~6_combout ;
wire \read_capture_delay_reg~12_combout ;
wire \read_capture_delay_reg[12]~q ;
wire \read_capture_delay_reg~11_combout ;
wire \read_capture_delay_reg[13]~q ;
wire \Mux0~7_combout ;
wire \read_capture_delay_reg~13_combout ;
wire \read_capture_delay_reg[14]~q ;
wire \Mux0~8_combout ;
wire \Mux0~9_combout ;
wire \Equal16~0_combout ;
wire \read_data_cnt~2_combout ;
wire \read_data_cnt~4_combout ;
wire \read_data_cnt[0]~1_combout ;
wire \read_data_cnt[0]~q ;
wire \Add6~1_combout ;
wire \read_data_cnt~3_combout ;
wire \read_data_cnt[1]~q ;
wire \Add6~0_combout ;
wire \read_data_cnt~0_combout ;
wire \read_data_cnt[2]~q ;
wire \read_data_done~0_combout ;
wire \read_data_cnt~5_combout ;
wire \read_data_cnt[3]~q ;
wire \read_data_done~combout ;
wire \read_data_valid~q ;
wire \flash_datain_reg~4_combout ;
wire \flash_datain_reg[0]~q ;
wire \flash_datain_reg~5_combout ;
wire \flash_datain_reg[1]~q ;
wire \Equal17~0_combout ;
wire \flash_datain_reg~6_combout ;
wire \flash_datain_reg[2]~q ;
wire \flash_datain_reg~7_combout ;
wire \flash_datain_reg[3]~q ;
wire \flash_datain_reg[4]~0_combout ;
wire \flash_datain_reg[4]~q ;
wire \flash_datain_reg[5]~1_combout ;
wire \flash_datain_reg[5]~q ;
wire \flash_datain_reg[6]~2_combout ;
wire \flash_datain_reg[6]~q ;
wire \flash_datain_reg[7]~3_combout ;
wire \flash_datain_reg[7]~q ;


flashLoader_clk_div clk_div_new_inst_2(
	.csr_clk_baud_rate_data_0(csr_clk_baud_rate_data_0),
	.reset(altera_reset_synchronizer_int_chain_out),
	.csr_clk_baud_rate_data_1(csr_clk_baud_rate_data_1),
	.csr_clk_baud_rate_data_2(csr_clk_baud_rate_data_2),
	.csr_clk_baud_rate_data_3(csr_clk_baud_rate_data_3),
	.csr_clk_baud_rate_data_4(csr_clk_baud_rate_data_4),
	.stateST_DEASSERT_CS_DLY(\state.ST_DEASSERT_CS_DLY~q ),
	.WideOr7(\WideOr7~0_combout ),
	.clk_track1(\clk_div_new_inst_2|clk_track~q ),
	.clk_out(\clk_div_new_inst_2|clk_out~0_combout ),
	.Equal0(\clk_div_new_inst_2|Equal0~1_combout ),
	.Equal01(\clk_div_new_inst_2|Equal0~2_combout ),
	.enable_d1(\clk_div_new_inst_2|enable_d~q ),
	.Add1(\clk_div_new_inst_2|Add1~1_combout ),
	.enable(\WideOr7~combout ),
	.Equal02(\clk_div_new_inst_2|Equal0~3_combout ),
	.rising_edge1(\clk_div_new_inst_2|rising_edge~combout ),
	.clk(clk_clk));

flashLoader_inf_sc_fifo_ser_data inf_sc_fifo_ser_data_inst(
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.out_payload_12(\inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|out_payload[12]~q ),
	.out_payload_2(\inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|out_payload[2]~q ),
	.out_payload_1(\inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|out_payload[1]~q ),
	.out_payload_0(\inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|out_payload[0]~q ),
	.mem_used_9(\inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|mem_used[9]~q ),
	.out_valid(\inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|out_valid~q ),
	.stateST_SEND(\state.ST_SEND~q ),
	.fifo_pop_out(\fifo_pop_out~1_combout ),
	.out_payload_16(\inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|out_payload[16]~q ),
	.out_payload_8(\inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|out_payload[8]~q ),
	.WideOr1(\qspi_inf_mux_inst|qspi_inf_mux|WideOr1~2_combout ),
	.write(\inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|write~0_combout ),
	.src_payload_0(\qspi_inf_mux_inst|qspi_inf_mux|src_payload[0]~1_combout ),
	.src_data_0(\qspi_inf_mux_inst|qspi_inf_mux|src_data[0]~1_combout ),
	.src_channel_2(\qspi_inf_mux_inst|qspi_inf_mux|src_channel[2]~1_combout ),
	.src_channel_1(\qspi_inf_mux_inst|qspi_inf_mux|src_channel[1]~3_combout ),
	.src_channel_0(\qspi_inf_mux_inst|qspi_inf_mux|src_channel[0]~5_combout ),
	.src_channel_8(\qspi_inf_mux_inst|qspi_inf_mux|src_channel[8]~7_combout ),
	.clk_clk(clk_clk));

flashLoader_qspi_inf_mux qspi_inf_mux_inst(
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.out_valid(\adapter_8_4_inst|out_valid~q ),
	.grant_0(\qspi_inf_mux_inst|qspi_inf_mux|arb|grant[0]~2_combout ),
	.out_valid1(\adapter_8_1_inst|out_valid~q ),
	.out_valid2(\adapter_8_2_inst|out_valid~q ),
	.request_1(\qspi_inf_mux_inst|qspi_inf_mux|request[1]~combout ),
	.full_addercout_1(\qspi_inf_mux_inst|qspi_inf_mux|arb|adder|full_adder.cout[1]~combout ),
	.cout(\qspi_inf_mux_inst|qspi_inf_mux|arb|adder|cout~0_combout ),
	.sum_1(\qspi_inf_mux_inst|qspi_inf_mux|arb|adder|sum[1]~combout ),
	.request_2(\qspi_inf_mux_inst|qspi_inf_mux|request[2]~combout ),
	.cout1(\qspi_inf_mux_inst|qspi_inf_mux|arb|adder|cout~1_combout ),
	.grant_01(\qspi_inf_mux_inst|qspi_inf_mux|arb|grant[0]~3_combout ),
	.WideOr1(\qspi_inf_mux_inst|qspi_inf_mux|WideOr1~2_combout ),
	.write(\inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|write~0_combout ),
	.out_endofpacket(\adapter_8_4_inst|out_endofpacket~q ),
	.out_endofpacket1(\adapter_8_1_inst|out_endofpacket~q ),
	.out_endofpacket2(\adapter_8_2_inst|out_endofpacket~q ),
	.src_payload_0(\qspi_inf_mux_inst|qspi_inf_mux|src_payload[0]~1_combout ),
	.out_data_0(\adapter_8_4_inst|out_data[0]~q ),
	.out_data_01(\adapter_8_1_inst|out_data[0]~q ),
	.out_data_02(\adapter_8_2_inst|out_data[0]~q ),
	.src_data_0(\qspi_inf_mux_inst|qspi_inf_mux|src_data[0]~1_combout ),
	.out_channel_2(\adapter_8_4_inst|out_channel[2]~q ),
	.out_channel_21(\adapter_8_1_inst|out_channel[2]~q ),
	.out_channel_22(\adapter_8_2_inst|out_channel[2]~q ),
	.src_channel_2(\qspi_inf_mux_inst|qspi_inf_mux|src_channel[2]~1_combout ),
	.out_channel_1(\adapter_8_4_inst|out_channel[1]~q ),
	.out_channel_11(\adapter_8_1_inst|out_channel[1]~q ),
	.out_channel_12(\adapter_8_2_inst|out_channel[1]~q ),
	.src_channel_1(\qspi_inf_mux_inst|qspi_inf_mux|src_channel[1]~3_combout ),
	.out_channel_0(\adapter_8_4_inst|out_channel[0]~q ),
	.out_channel_01(\adapter_8_1_inst|out_channel[0]~q ),
	.out_channel_02(\adapter_8_2_inst|out_channel[0]~q ),
	.src_channel_0(\qspi_inf_mux_inst|qspi_inf_mux|src_channel[0]~5_combout ),
	.out_channel_8(\adapter_8_4_inst|out_channel[8]~q ),
	.out_channel_81(\adapter_8_1_inst|out_channel[8]~q ),
	.out_channel_82(\adapter_8_2_inst|out_channel[8]~q ),
	.src_channel_8(\qspi_inf_mux_inst|qspi_inf_mux|src_channel[8]~7_combout ),
	.clk_clk(clk_clk));

flashLoader_adapter_8_4 adapter_8_4_inst(
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.in_channel({gnd,gnd,gnd,Selector17,gnd,gnd,gnd,gnd,gnd,stateST_SEND_DATA,stateST_SEND_ADDR,stateST_SEND_OPCODE}),
	.out_valid1(\adapter_8_4_inst|out_valid~q ),
	.request_1(\qspi_inf_mux_inst|qspi_inf_mux|request[1]~combout ),
	.full_addercout_1(\qspi_inf_mux_inst|qspi_inf_mux|arb|adder|full_adder.cout[1]~combout ),
	.cout(\qspi_inf_mux_inst|qspi_inf_mux|arb|adder|cout~0_combout ),
	.mem_used_9(\inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|mem_used[9]~q ),
	.request_2(\qspi_inf_mux_inst|qspi_inf_mux|request[2]~combout ),
	.cout1(\qspi_inf_mux_inst|qspi_inf_mux|arb|adder|cout~1_combout ),
	.state_register_0(\adapter_8_4_inst|state_register[0]~q ),
	.always4(\adapter_8_4_inst|always4~0_combout ),
	.always41(\adapter_8_4_inst|always4~1_combout ),
	.a_valid1(\adapter_8_4_inst|a_valid~q ),
	.in_ready1(in_ready),
	.out_endofpacket1(\adapter_8_4_inst|out_endofpacket~q ),
	.in_valid(\demultiplexer_inst|src2_valid~combout ),
	.out_data_0(\adapter_8_4_inst|out_data[0]~q ),
	.out_channel_2(\adapter_8_4_inst|out_channel[2]~q ),
	.out_channel_1(\adapter_8_4_inst|out_channel[1]~q ),
	.out_channel_0(\adapter_8_4_inst|out_channel[0]~q ),
	.out_channel_8(\adapter_8_4_inst|out_channel[8]~q ),
	.in_endofpacket(Selector20),
	.in_data({gnd,gnd,gnd,Selector12,gnd,gnd,gnd,Selector16}),
	.clk(clk_clk));

flashLoader_adapter_8_2 adapter_8_2_inst(
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.in_channel({gnd,gnd,gnd,Selector17,gnd,gnd,gnd,gnd,gnd,stateST_SEND_DATA,stateST_SEND_ADDR,stateST_SEND_OPCODE}),
	.out_valid1(\adapter_8_2_inst|out_valid~q ),
	.request_1(\qspi_inf_mux_inst|qspi_inf_mux|request[1]~combout ),
	.mem_used_9(\inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|mem_used[9]~q ),
	.state_register_1(\adapter_8_2_inst|state_register[1]~q ),
	.state_register_0(\adapter_8_2_inst|state_register[0]~q ),
	.a_valid1(\adapter_8_2_inst|a_valid~q ),
	.sum_1(\qspi_inf_mux_inst|qspi_inf_mux|arb|adder|sum[1]~combout ),
	.cout(\qspi_inf_mux_inst|qspi_inf_mux|arb|adder|cout~1_combout ),
	.always4(\adapter_8_2_inst|always4~1_combout ),
	.in_ready1(\adapter_8_2_inst|in_ready~combout ),
	.out_endofpacket1(\adapter_8_2_inst|out_endofpacket~q ),
	.in_valid(\demultiplexer_inst|src1_valid~combout ),
	.out_data_0(\adapter_8_2_inst|out_data[0]~q ),
	.out_channel_2(\adapter_8_2_inst|out_channel[2]~q ),
	.out_channel_1(\adapter_8_2_inst|out_channel[1]~q ),
	.out_channel_0(\adapter_8_2_inst|out_channel[0]~q ),
	.out_channel_8(\adapter_8_2_inst|out_channel[8]~q ),
	.in_endofpacket(Selector20),
	.in_data({gnd,Selector10,gnd,Selector12,gnd,Selector14,gnd,Selector16}),
	.clk(clk_clk));

flashLoader_adapter_8_1 adapter_8_1_inst(
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.in_channel({gnd,gnd,gnd,Selector17,gnd,gnd,gnd,gnd,gnd,stateST_SEND_DATA,stateST_SEND_ADDR,stateST_SEND_OPCODE}),
	.grant_0(\qspi_inf_mux_inst|qspi_inf_mux|arb|grant[0]~2_combout ),
	.out_valid1(\adapter_8_1_inst|out_valid~q ),
	.full_addercout_1(\qspi_inf_mux_inst|qspi_inf_mux|arb|adder|full_adder.cout[1]~combout ),
	.cout(\qspi_inf_mux_inst|qspi_inf_mux|arb|adder|cout~0_combout ),
	.mem_used_9(\inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|mem_used[9]~q ),
	.in_ready1(\adapter_8_1_inst|in_ready~combout ),
	.grant_01(\qspi_inf_mux_inst|qspi_inf_mux|arb|grant[0]~3_combout ),
	.out_endofpacket1(\adapter_8_1_inst|out_endofpacket~q ),
	.in_valid(\demultiplexer_inst|src0_valid~combout ),
	.out_data_0(\adapter_8_1_inst|out_data[0]~q ),
	.out_channel_2(\adapter_8_1_inst|out_channel[2]~q ),
	.out_channel_1(\adapter_8_1_inst|out_channel[1]~q ),
	.out_channel_0(\adapter_8_1_inst|out_channel[0]~q ),
	.out_channel_8(\adapter_8_1_inst|out_channel[8]~q ),
	.in_endofpacket(Selector20),
	.in_data({Selector9,Selector10,Selector11,Selector12,Selector13,Selector14,Selector15,Selector16}),
	.clk(clk_clk));

flashLoader_demultiplexer_12_channels demultiplexer_inst(
	.data_num_lines_1(data_num_lines_1),
	.data_num_lines_2(data_num_lines_2),
	.addr_num_lines_2(addr_num_lines_2),
	.addr_num_lines_1(addr_num_lines_1),
	.in_cmd_channel_reg_1(in_cmd_channel_reg_1),
	.in_cmd_channel_reg_0(in_cmd_channel_reg_0),
	.op_num_lines_1(op_num_lines_1),
	.in_ready(\adapter_8_1_inst|in_ready~combout ),
	.data_num_lines_0(data_num_lines_0),
	.op_num_lines_0(op_num_lines_0),
	.state_register_1(\adapter_8_2_inst|state_register[1]~q ),
	.state_register_0(\adapter_8_2_inst|state_register[0]~q ),
	.a_valid(\adapter_8_2_inst|a_valid~q ),
	.always4(\adapter_8_2_inst|always4~1_combout ),
	.WideOr0(WideOr0),
	.state_register_01(\adapter_8_4_inst|state_register[0]~q ),
	.always41(\adapter_8_4_inst|always4~0_combout ),
	.always42(\adapter_8_4_inst|always4~1_combout ),
	.a_valid1(\adapter_8_4_inst|a_valid~q ),
	.in_ready1(in_ready),
	.op_num_lines_2(op_num_lines_2),
	.WideOr01(WideOr01),
	.Selector8(Selector8),
	.demux_channel_2(\demux_channel[2]~0_combout ),
	.Equal0(\Equal0~0_combout ),
	.demux_channel_21(demux_channel_2),
	.sink_ready(in_cmd_ready),
	.in_ready2(\adapter_8_2_inst|in_ready~combout ),
	.demux_channel_1(\demux_channel[1]~2_combout ),
	.demux_channel_11(\demux_channel[1]~3_combout ),
	.addr_num_lines_0(addr_num_lines_0),
	.demux_channel_0(\demux_channel[0]~4_combout ),
	.demux_channel_01(\demux_channel[0]~5_combout ),
	.WideOr02(WideOr02),
	.WideOr03(WideOr03),
	.WideOr04(WideOr04),
	.WideOr05(WideOr05),
	.demux_channel_22(\demux_channel[2]~6_combout ),
	.src0_valid1(\demultiplexer_inst|src0_valid~combout ),
	.src1_valid1(\demultiplexer_inst|src1_valid~combout ),
	.src2_valid1(\demultiplexer_inst|src2_valid~combout ),
	.WideOr06(WideOr06));

cycloneive_lcell_comb \WideOr7~0 (
	.dataa(\state.ST_DEASSERT_CS~q ),
	.datab(\state.ST_ASSERT_CS_DLY~q ),
	.datac(\state.ST_STOP_CLK~q ),
	.datad(\state.ST_IDLE~q ),
	.cin(gnd),
	.combout(\WideOr7~0_combout ),
	.cout());
defparam \WideOr7~0 .lut_mask = 16'hFEFF;
defparam \WideOr7~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb WideOr7(
	.dataa(\state.ST_DEASSERT_CS_DLY~q ),
	.datab(\WideOr7~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\WideOr7~combout ),
	.cout());
defparam WideOr7.lut_mask = 16'h1111;
defparam WideOr7.sum_lutc_input = "datac";

cycloneive_lcell_comb \demux_channel[1]~2 (
	.dataa(addr_num_lines_1),
	.datab(data_num_lines_1),
	.datac(gnd),
	.datad(stateST_SEND_ADDR),
	.cin(gnd),
	.combout(\demux_channel[1]~2_combout ),
	.cout());
defparam \demux_channel[1]~2 .lut_mask = 16'hAACC;
defparam \demux_channel[1]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \demux_channel[1]~3 (
	.dataa(op_num_lines_1),
	.datab(\demux_channel[1]~2_combout ),
	.datac(\Equal0~0_combout ),
	.datad(stateST_SEND_OPCODE),
	.cin(gnd),
	.combout(\demux_channel[1]~3_combout ),
	.cout());
defparam \demux_channel[1]~3 .lut_mask = 16'hAAAC;
defparam \demux_channel[1]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \demux_channel[0]~4 (
	.dataa(addr_num_lines_0),
	.datab(data_num_lines_0),
	.datac(gnd),
	.datad(stateST_SEND_ADDR),
	.cin(gnd),
	.combout(\demux_channel[0]~4_combout ),
	.cout());
defparam \demux_channel[0]~4 .lut_mask = 16'hAACC;
defparam \demux_channel[0]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \demux_channel[0]~5 (
	.dataa(op_num_lines_0),
	.datab(\demux_channel[0]~4_combout ),
	.datac(\Equal0~0_combout ),
	.datad(stateST_SEND_OPCODE),
	.cin(gnd),
	.combout(\demux_channel[0]~5_combout ),
	.cout());
defparam \demux_channel[0]~5 .lut_mask = 16'hAAAC;
defparam \demux_channel[0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \demux_channel[2]~6 (
	.dataa(stateST_SEND_OPCODE),
	.datab(in_cmd_channel_reg_1),
	.datac(gnd),
	.datad(in_cmd_channel_reg_0),
	.cin(gnd),
	.combout(\demux_channel[2]~6_combout ),
	.cout());
defparam \demux_channel[2]~6 .lut_mask = 16'hAAEE;
defparam \demux_channel[2]~6 .sum_lutc_input = "datac";

dffeas flash_clk_reg(
	.clk(clk_clk),
	.d(\clk_div_new_inst_2|clk_out~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(flash_clk_reg1),
	.prn(vcc));
defparam flash_clk_reg.is_wysiwyg = "true";
defparam flash_clk_reg.power_up = "low";

dffeas oe_reg(
	.clk(clk_clk),
	.d(qspi_interface_en),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oe_reg1),
	.prn(vcc));
defparam oe_reg.is_wysiwyg = "true";
defparam oe_reg.power_up = "low";

dffeas \ncs_reg[0] (
	.clk(clk_clk),
	.d(\ncs_wire[0]~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ncs_reg_0),
	.prn(vcc));
defparam \ncs_reg[0] .is_wysiwyg = "true";
defparam \ncs_reg[0] .power_up = "low";

dffeas \flash_data_out_reg[0] (
	.clk(clk_clk),
	.d(\flash_data_out[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(flash_data_out_reg_0),
	.prn(vcc));
defparam \flash_data_out_reg[0] .is_wysiwyg = "true";
defparam \flash_data_out_reg[0] .power_up = "low";

cycloneive_lcell_comb \demux_channel[2]~1 (
	.dataa(op_num_lines_2),
	.datab(\demux_channel[2]~0_combout ),
	.datac(\Equal0~0_combout ),
	.datad(stateST_SEND_OPCODE),
	.cin(gnd),
	.combout(demux_channel_2),
	.cout());
defparam \demux_channel[2]~1 .lut_mask = 16'hAAAC;
defparam \demux_channel[2]~1 .sum_lutc_input = "datac";

dffeas out_rsp_valid(
	.clk(clk_clk),
	.d(\read_data_valid~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_rsp_valid1),
	.prn(vcc));
defparam out_rsp_valid.is_wysiwyg = "true";
defparam out_rsp_valid.power_up = "low";

dffeas \out_rsp_data[0] (
	.clk(clk_clk),
	.d(\flash_datain_reg[0]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_valid~q ),
	.q(out_rsp_data_0),
	.prn(vcc));
defparam \out_rsp_data[0] .is_wysiwyg = "true";
defparam \out_rsp_data[0] .power_up = "low";

dffeas \out_rsp_data[1] (
	.clk(clk_clk),
	.d(\flash_datain_reg[1]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_valid~q ),
	.q(out_rsp_data_1),
	.prn(vcc));
defparam \out_rsp_data[1] .is_wysiwyg = "true";
defparam \out_rsp_data[1] .power_up = "low";

dffeas \out_rsp_data[2] (
	.clk(clk_clk),
	.d(\flash_datain_reg[2]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_valid~q ),
	.q(out_rsp_data_2),
	.prn(vcc));
defparam \out_rsp_data[2] .is_wysiwyg = "true";
defparam \out_rsp_data[2] .power_up = "low";

dffeas \out_rsp_data[3] (
	.clk(clk_clk),
	.d(\flash_datain_reg[3]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_valid~q ),
	.q(out_rsp_data_3),
	.prn(vcc));
defparam \out_rsp_data[3] .is_wysiwyg = "true";
defparam \out_rsp_data[3] .power_up = "low";

dffeas \out_rsp_data[4] (
	.clk(clk_clk),
	.d(\flash_datain_reg[4]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_valid~q ),
	.q(out_rsp_data_4),
	.prn(vcc));
defparam \out_rsp_data[4] .is_wysiwyg = "true";
defparam \out_rsp_data[4] .power_up = "low";

dffeas \out_rsp_data[5] (
	.clk(clk_clk),
	.d(\flash_datain_reg[5]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_valid~q ),
	.q(out_rsp_data_5),
	.prn(vcc));
defparam \out_rsp_data[5] .is_wysiwyg = "true";
defparam \out_rsp_data[5] .power_up = "low";

dffeas \out_rsp_data[6] (
	.clk(clk_clk),
	.d(\flash_datain_reg[6]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_valid~q ),
	.q(out_rsp_data_6),
	.prn(vcc));
defparam \out_rsp_data[6] .is_wysiwyg = "true";
defparam \out_rsp_data[6] .power_up = "low";

dffeas \out_rsp_data[7] (
	.clk(clk_clk),
	.d(\flash_datain_reg[7]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_valid~q ),
	.q(out_rsp_data_7),
	.prn(vcc));
defparam \out_rsp_data[7] .is_wysiwyg = "true";
defparam \out_rsp_data[7] .power_up = "low";

cycloneive_lcell_comb \Selector0~0 (
	.dataa(\state.ST_DEASSERT_CS~q ),
	.datab(gnd),
	.datac(\state.ST_IDLE~q ),
	.datad(\inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|out_valid~q ),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
defparam \Selector0~0 .lut_mask = 16'h5550;
defparam \Selector0~0 .sum_lutc_input = "datac";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_IDLE~q ),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cycloneive_lcell_comb \LessThan0~0 (
	.dataa(\inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|out_valid~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\state.ST_IDLE~q ),
	.cin(gnd),
	.combout(\LessThan0~0_combout ),
	.cout());
defparam \LessThan0~0 .lut_mask = 16'h00AA;
defparam \LessThan0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal14~1 (
	.dataa(csr_delay_setting_data_1),
	.datab(csr_delay_setting_data_2),
	.datac(\cs_assert_cnt[2]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal14~1_combout ),
	.cout());
defparam \Equal14~1 .lut_mask = 16'h9696;
defparam \Equal14~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cs_assert_cnt_next~4 (
	.dataa(gnd),
	.datab(\cs_assert_cnt[0]~q ),
	.datac(\cs_assert_cnt[1]~q ),
	.datad(\Equal14~3_combout ),
	.cin(gnd),
	.combout(\cs_assert_cnt_next~4_combout ),
	.cout());
defparam \cs_assert_cnt_next~4 .lut_mask = 16'h003C;
defparam \cs_assert_cnt_next~4 .sum_lutc_input = "datac";

dffeas \cs_assert_cnt[1] (
	.clk(clk_clk),
	.d(\cs_assert_cnt_next~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.ST_ASSERT_CS_DLY~q ),
	.q(\cs_assert_cnt[1]~q ),
	.prn(vcc));
defparam \cs_assert_cnt[1] .is_wysiwyg = "true";
defparam \cs_assert_cnt[1] .power_up = "low";

cycloneive_lcell_comb \Equal14~2 (
	.dataa(csr_delay_setting_data_0),
	.datab(\cs_assert_cnt[0]~q ),
	.datac(csr_delay_setting_data_1),
	.datad(\cs_assert_cnt[1]~q ),
	.cin(gnd),
	.combout(\Equal14~2_combout ),
	.cout());
defparam \Equal14~2 .lut_mask = 16'h0990;
defparam \Equal14~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cs_assert_cnt_next~3 (
	.dataa(\cs_assert_cnt[0]~q ),
	.datab(\Equal14~0_combout ),
	.datac(\Equal14~1_combout ),
	.datad(\Equal14~2_combout ),
	.cin(gnd),
	.combout(\cs_assert_cnt_next~3_combout ),
	.cout());
defparam \cs_assert_cnt_next~3 .lut_mask = 16'h1555;
defparam \cs_assert_cnt_next~3 .sum_lutc_input = "datac";

dffeas \cs_assert_cnt[0] (
	.clk(clk_clk),
	.d(\cs_assert_cnt_next~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.ST_ASSERT_CS_DLY~q ),
	.q(\cs_assert_cnt[0]~q ),
	.prn(vcc));
defparam \cs_assert_cnt[0] .is_wysiwyg = "true";
defparam \cs_assert_cnt[0] .power_up = "low";

cycloneive_lcell_comb \cs_assert_cnt_next~5 (
	.dataa(\cs_assert_cnt[0]~q ),
	.datab(\cs_assert_cnt[1]~q ),
	.datac(\cs_assert_cnt[2]~q ),
	.datad(\Equal14~3_combout ),
	.cin(gnd),
	.combout(\cs_assert_cnt_next~5_combout ),
	.cout());
defparam \cs_assert_cnt_next~5 .lut_mask = 16'h0078;
defparam \cs_assert_cnt_next~5 .sum_lutc_input = "datac";

dffeas \cs_assert_cnt[2] (
	.clk(clk_clk),
	.d(\cs_assert_cnt_next~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.ST_ASSERT_CS_DLY~q ),
	.q(\cs_assert_cnt[2]~q ),
	.prn(vcc));
defparam \cs_assert_cnt[2] .is_wysiwyg = "true";
defparam \cs_assert_cnt[2] .power_up = "low";

cycloneive_lcell_comb \Add3~0 (
	.dataa(\cs_assert_cnt[0]~q ),
	.datab(\cs_assert_cnt[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add3~0_combout ),
	.cout());
defparam \Add3~0 .lut_mask = 16'h8888;
defparam \Add3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cs_assert_cnt_next~2 (
	.dataa(\cs_assert_cnt[3]~q ),
	.datab(\cs_assert_cnt[2]~q ),
	.datac(\Add3~0_combout ),
	.datad(\Equal14~3_combout ),
	.cin(gnd),
	.combout(\cs_assert_cnt_next~2_combout ),
	.cout());
defparam \cs_assert_cnt_next~2 .lut_mask = 16'h006A;
defparam \cs_assert_cnt_next~2 .sum_lutc_input = "datac";

dffeas \cs_assert_cnt[3] (
	.clk(clk_clk),
	.d(\cs_assert_cnt_next~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.ST_ASSERT_CS_DLY~q ),
	.q(\cs_assert_cnt[3]~q ),
	.prn(vcc));
defparam \cs_assert_cnt[3] .is_wysiwyg = "true";
defparam \cs_assert_cnt[3] .power_up = "low";

cycloneive_lcell_comb \Equal14~0 (
	.dataa(csr_delay_setting_data_3),
	.datab(\cs_assert_cnt[3]~q ),
	.datac(csr_delay_setting_data_1),
	.datad(csr_delay_setting_data_2),
	.cin(gnd),
	.combout(\Equal14~0_combout ),
	.cout());
defparam \Equal14~0 .lut_mask = 16'h9996;
defparam \Equal14~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal14~3 (
	.dataa(\Equal14~0_combout ),
	.datab(\Equal14~1_combout ),
	.datac(\Equal14~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal14~3_combout ),
	.cout());
defparam \Equal14~3 .lut_mask = 16'h8080;
defparam \Equal14~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ncs_wire[0]~2 (
	.dataa(gnd),
	.datab(csr_delay_setting_data_1),
	.datac(csr_delay_setting_data_2),
	.datad(csr_delay_setting_data_3),
	.cin(gnd),
	.combout(\ncs_wire[0]~2_combout ),
	.cout());
defparam \ncs_wire[0]~2 .lut_mask = 16'h0003;
defparam \ncs_wire[0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~0 (
	.dataa(\state.ST_ASSERT_CS_DLY~q ),
	.datab(\LessThan0~0_combout ),
	.datac(\Equal14~3_combout ),
	.datad(\ncs_wire[0]~2_combout ),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'h0ACE;
defparam \Selector1~0 .sum_lutc_input = "datac";

dffeas \state.ST_ASSERT_CS_DLY (
	.clk(clk_clk),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_ASSERT_CS_DLY~q ),
	.prn(vcc));
defparam \state.ST_ASSERT_CS_DLY .is_wysiwyg = "true";
defparam \state.ST_ASSERT_CS_DLY .power_up = "low";

cycloneive_lcell_comb \Selector2~0 (
	.dataa(\state.ST_ASSERT_CS_DLY~q ),
	.datab(\ncs_wire[0]~2_combout ),
	.datac(\LessThan0~0_combout ),
	.datad(\Equal14~3_combout ),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
defparam \Selector2~0 .lut_mask = 16'hEAC0;
defparam \Selector2~0 .sum_lutc_input = "datac";

dffeas \state.ST_START_CLK (
	.clk(clk_clk),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_START_CLK~q ),
	.prn(vcc));
defparam \state.ST_START_CLK .is_wysiwyg = "true";
defparam \state.ST_START_CLK .power_up = "low";

cycloneive_lcell_comb \require_rdata_reg~0 (
	.dataa(stateST_IDLE),
	.datab(header_information_11),
	.datac(\require_rdata_reg~q ),
	.datad(\state.ST_START_CLK~q ),
	.cin(gnd),
	.combout(\require_rdata_reg~0_combout ),
	.cout());
defparam \require_rdata_reg~0 .lut_mask = 16'h88F0;
defparam \require_rdata_reg~0 .sum_lutc_input = "datac";

dffeas require_rdata_reg(
	.clk(clk_clk),
	.d(\require_rdata_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\require_rdata_reg~q ),
	.prn(vcc));
defparam require_rdata_reg.is_wysiwyg = "true";
defparam require_rdata_reg.power_up = "low";

dffeas \state.ST_ASSERT_CS (
	.clk(clk_clk),
	.d(\state.ST_START_CLK~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_ASSERT_CS~q ),
	.prn(vcc));
defparam \state.ST_ASSERT_CS .is_wysiwyg = "true";
defparam \state.ST_ASSERT_CS .power_up = "low";

cycloneive_lcell_comb \fifo_pop_out~0 (
	.dataa(\clk_div_new_inst_2|enable_d~q ),
	.datab(csr_clk_baud_rate_data_3),
	.datac(\clk_div_new_inst_2|Add1~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\fifo_pop_out~0_combout ),
	.cout());
defparam \fifo_pop_out~0 .lut_mask = 16'h8282;
defparam \fifo_pop_out~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_pop_out~1 (
	.dataa(\clk_div_new_inst_2|clk_track~q ),
	.datab(\clk_div_new_inst_2|Equal0~1_combout ),
	.datac(\clk_div_new_inst_2|Equal0~2_combout ),
	.datad(\fifo_pop_out~0_combout ),
	.cin(gnd),
	.combout(\fifo_pop_out~1_combout ),
	.cout());
defparam \fifo_pop_out~1 .lut_mask = 16'h4000;
defparam \fifo_pop_out~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_state~1 (
	.dataa(\inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|out_payload[16]~q ),
	.datab(\inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|out_payload[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_state~1_combout ),
	.cout());
defparam \next_state~1 .lut_mask = 16'h8888;
defparam \next_state~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector3~0 (
	.dataa(\state.ST_ASSERT_CS~q ),
	.datab(\state.ST_SEND~q ),
	.datac(\fifo_pop_out~1_combout ),
	.datad(\next_state~1_combout ),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
defparam \Selector3~0 .lut_mask = 16'hAEEE;
defparam \Selector3~0 .sum_lutc_input = "datac";

dffeas \state.ST_SEND (
	.clk(clk_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_SEND~q ),
	.prn(vcc));
defparam \state.ST_SEND .is_wysiwyg = "true";
defparam \state.ST_SEND .power_up = "low";

cycloneive_lcell_comb \next_state~0 (
	.dataa(\state.ST_SEND~q ),
	.datab(\fifo_pop_out~1_combout ),
	.datac(\inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|out_payload[16]~q ),
	.datad(\inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|out_payload[8]~q ),
	.cin(gnd),
	.combout(\next_state~0_combout ),
	.cout());
defparam \next_state~0 .lut_mask = 16'h8000;
defparam \next_state~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \LessThan1~0 (
	.dataa(header_information_17),
	.datab(header_information_16),
	.datac(header_information_15),
	.datad(header_information_14),
	.cin(gnd),
	.combout(\LessThan1~0_combout ),
	.cout());
defparam \LessThan1~0 .lut_mask = 16'hFFFE;
defparam \LessThan1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector5~0 (
	.dataa(\require_rdata_reg~q ),
	.datab(\next_state~0_combout ),
	.datac(header_information_13),
	.datad(\LessThan1~0_combout ),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
defparam \Selector5~0 .lut_mask = 16'h0008;
defparam \Selector5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector5~1 (
	.dataa(stateST_IDLE),
	.datab(\state.ST_RECEIVE~q ),
	.datac(header_information_11),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector5~1_combout ),
	.cout());
defparam \Selector5~1 .lut_mask = 16'h8080;
defparam \Selector5~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_state~2 (
	.dataa(\require_rdata_reg~q ),
	.datab(\next_state~0_combout ),
	.datac(header_information_13),
	.datad(\LessThan1~0_combout ),
	.cin(gnd),
	.combout(\next_state~2_combout ),
	.cout());
defparam \next_state~2 .lut_mask = 16'h8880;
defparam \next_state~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~0 (
	.dataa(header_information_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
defparam \Add0~0 .lut_mask = 16'h55AA;
defparam \Add0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~2 (
	.dataa(header_information_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
defparam \Add0~2 .lut_mask = 16'hA505;
defparam \Add0~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~4 (
	.dataa(header_information_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
defparam \Add0~4 .lut_mask = 16'h5AAF;
defparam \Add0~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~6 (
	.dataa(header_information_16),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
defparam \Add0~6 .lut_mask = 16'hA505;
defparam \Add0~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~8 (
	.dataa(header_information_17),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout());
defparam \Add0~8 .lut_mask = 16'h5A5A;
defparam \Add0~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \dummy_cnt[0]~5 (
	.dataa(\dummy_cnt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\dummy_cnt[0]~5_combout ),
	.cout(\dummy_cnt[0]~6 ));
defparam \dummy_cnt[0]~5 .lut_mask = 16'h55AA;
defparam \dummy_cnt[0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always6~1 (
	.dataa(\clk_div_new_inst_2|Equal0~3_combout ),
	.datab(\clk_div_new_inst_2|enable_d~q ),
	.datac(\state.ST_DUMMY_CYCLES~q ),
	.datad(\clk_div_new_inst_2|clk_track~q ),
	.cin(gnd),
	.combout(\always6~1_combout ),
	.cout());
defparam \always6~1 .lut_mask = 16'h0080;
defparam \always6~1 .sum_lutc_input = "datac";

dffeas \dummy_cnt[0] (
	.clk(clk_clk),
	.d(\dummy_cnt[0]~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(\dummy_cnt_done~3_combout ),
	.sload(gnd),
	.ena(\always6~1_combout ),
	.q(\dummy_cnt[0]~q ),
	.prn(vcc));
defparam \dummy_cnt[0] .is_wysiwyg = "true";
defparam \dummy_cnt[0] .power_up = "low";

cycloneive_lcell_comb \dummy_cnt[1]~7 (
	.dataa(\dummy_cnt[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\dummy_cnt[0]~6 ),
	.combout(\dummy_cnt[1]~7_combout ),
	.cout(\dummy_cnt[1]~8 ));
defparam \dummy_cnt[1]~7 .lut_mask = 16'h5A5F;
defparam \dummy_cnt[1]~7 .sum_lutc_input = "cin";

dffeas \dummy_cnt[1] (
	.clk(clk_clk),
	.d(\dummy_cnt[1]~7_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(\dummy_cnt_done~3_combout ),
	.sload(gnd),
	.ena(\always6~1_combout ),
	.q(\dummy_cnt[1]~q ),
	.prn(vcc));
defparam \dummy_cnt[1] .is_wysiwyg = "true";
defparam \dummy_cnt[1] .power_up = "low";

cycloneive_lcell_comb \dummy_cnt[2]~9 (
	.dataa(\dummy_cnt[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\dummy_cnt[1]~8 ),
	.combout(\dummy_cnt[2]~9_combout ),
	.cout(\dummy_cnt[2]~10 ));
defparam \dummy_cnt[2]~9 .lut_mask = 16'hA50A;
defparam \dummy_cnt[2]~9 .sum_lutc_input = "cin";

dffeas \dummy_cnt[2] (
	.clk(clk_clk),
	.d(\dummy_cnt[2]~9_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(\dummy_cnt_done~3_combout ),
	.sload(gnd),
	.ena(\always6~1_combout ),
	.q(\dummy_cnt[2]~q ),
	.prn(vcc));
defparam \dummy_cnt[2] .is_wysiwyg = "true";
defparam \dummy_cnt[2] .power_up = "low";

cycloneive_lcell_comb \dummy_cnt[3]~11 (
	.dataa(\dummy_cnt[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\dummy_cnt[2]~10 ),
	.combout(\dummy_cnt[3]~11_combout ),
	.cout(\dummy_cnt[3]~12 ));
defparam \dummy_cnt[3]~11 .lut_mask = 16'h5A5F;
defparam \dummy_cnt[3]~11 .sum_lutc_input = "cin";

dffeas \dummy_cnt[3] (
	.clk(clk_clk),
	.d(\dummy_cnt[3]~11_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(\dummy_cnt_done~3_combout ),
	.sload(gnd),
	.ena(\always6~1_combout ),
	.q(\dummy_cnt[3]~q ),
	.prn(vcc));
defparam \dummy_cnt[3] .is_wysiwyg = "true";
defparam \dummy_cnt[3] .power_up = "low";

cycloneive_lcell_comb \dummy_cnt[4]~13 (
	.dataa(\dummy_cnt[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\dummy_cnt[3]~12 ),
	.combout(\dummy_cnt[4]~13_combout ),
	.cout());
defparam \dummy_cnt[4]~13 .lut_mask = 16'hA5A5;
defparam \dummy_cnt[4]~13 .sum_lutc_input = "cin";

dffeas \dummy_cnt[4] (
	.clk(clk_clk),
	.d(\dummy_cnt[4]~13_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(\dummy_cnt_done~3_combout ),
	.sload(gnd),
	.ena(\always6~1_combout ),
	.q(\dummy_cnt[4]~q ),
	.prn(vcc));
defparam \dummy_cnt[4] .is_wysiwyg = "true";
defparam \dummy_cnt[4] .power_up = "low";

cycloneive_lcell_comb \dummy_cnt_done~0 (
	.dataa(\Add0~4_combout ),
	.datab(\Add0~6_combout ),
	.datac(\dummy_cnt[3]~q ),
	.datad(\dummy_cnt[2]~q ),
	.cin(gnd),
	.combout(\dummy_cnt_done~0_combout ),
	.cout());
defparam \dummy_cnt_done~0 .lut_mask = 16'h8241;
defparam \dummy_cnt_done~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \dummy_cnt_done~1 (
	.dataa(\Add0~0_combout ),
	.datab(\Add0~2_combout ),
	.datac(\dummy_cnt[1]~q ),
	.datad(\dummy_cnt[0]~q ),
	.cin(gnd),
	.combout(\dummy_cnt_done~1_combout ),
	.cout());
defparam \dummy_cnt_done~1 .lut_mask = 16'h8241;
defparam \dummy_cnt_done~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \dummy_cnt_done~2 (
	.dataa(\fifo_pop_out~1_combout ),
	.datab(\dummy_cnt_done~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\dummy_cnt_done~2_combout ),
	.cout());
defparam \dummy_cnt_done~2 .lut_mask = 16'h8888;
defparam \dummy_cnt_done~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \dummy_cnt_done~3 (
	.dataa(\Add0~8_combout ),
	.datab(\dummy_cnt[4]~q ),
	.datac(\dummy_cnt_done~0_combout ),
	.datad(\dummy_cnt_done~2_combout ),
	.cin(gnd),
	.combout(\dummy_cnt_done~3_combout ),
	.cout());
defparam \dummy_cnt_done~3 .lut_mask = 16'h9000;
defparam \dummy_cnt_done~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector4~0 (
	.dataa(\next_state~2_combout ),
	.datab(\state.ST_DUMMY_CYCLES~q ),
	.datac(gnd),
	.datad(\dummy_cnt_done~3_combout ),
	.cin(gnd),
	.combout(\Selector4~0_combout ),
	.cout());
defparam \Selector4~0 .lut_mask = 16'hAAEE;
defparam \Selector4~0 .sum_lutc_input = "datac";

dffeas \state.ST_DUMMY_CYCLES (
	.clk(clk_clk),
	.d(\Selector4~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_DUMMY_CYCLES~q ),
	.prn(vcc));
defparam \state.ST_DUMMY_CYCLES .is_wysiwyg = "true";
defparam \state.ST_DUMMY_CYCLES .power_up = "low";

cycloneive_lcell_comb \Selector5~2 (
	.dataa(\Selector5~0_combout ),
	.datab(\Selector5~1_combout ),
	.datac(\state.ST_DUMMY_CYCLES~q ),
	.datad(\dummy_cnt_done~3_combout ),
	.cin(gnd),
	.combout(\Selector5~2_combout ),
	.cout());
defparam \Selector5~2 .lut_mask = 16'hFEEE;
defparam \Selector5~2 .sum_lutc_input = "datac";

dffeas \state.ST_RECEIVE (
	.clk(clk_clk),
	.d(\Selector5~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_RECEIVE~q ),
	.prn(vcc));
defparam \state.ST_RECEIVE .is_wysiwyg = "true";
defparam \state.ST_RECEIVE .power_up = "low";

cycloneive_lcell_comb \Selector6~0 (
	.dataa(\state.ST_RECEIVE~q ),
	.datab(gnd),
	.datac(stateST_IDLE),
	.datad(header_information_11),
	.cin(gnd),
	.combout(\Selector6~0_combout ),
	.cout());
defparam \Selector6~0 .lut_mask = 16'h0AAA;
defparam \Selector6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector6~1 (
	.dataa(\Selector6~0_combout ),
	.datab(\next_state~0_combout ),
	.datac(gnd),
	.datad(\require_rdata_reg~q ),
	.cin(gnd),
	.combout(\Selector6~1_combout ),
	.cout());
defparam \Selector6~1 .lut_mask = 16'hAAEE;
defparam \Selector6~1 .sum_lutc_input = "datac";

dffeas \state.ST_STOP_CLK (
	.clk(clk_clk),
	.d(\Selector6~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_STOP_CLK~q ),
	.prn(vcc));
defparam \state.ST_STOP_CLK .is_wysiwyg = "true";
defparam \state.ST_STOP_CLK .power_up = "low";

cycloneive_lcell_comb \cs_deassert_cnt_next~4 (
	.dataa(gnd),
	.datab(\cs_deassert_cnt[0]~q ),
	.datac(\cs_deassert_cnt[1]~q ),
	.datad(\Equal15~3_combout ),
	.cin(gnd),
	.combout(\cs_deassert_cnt_next~4_combout ),
	.cout());
defparam \cs_deassert_cnt_next~4 .lut_mask = 16'h003C;
defparam \cs_deassert_cnt_next~4 .sum_lutc_input = "datac";

dffeas \cs_deassert_cnt[1] (
	.clk(clk_clk),
	.d(\cs_deassert_cnt_next~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.ST_DEASSERT_CS_DLY~q ),
	.q(\cs_deassert_cnt[1]~q ),
	.prn(vcc));
defparam \cs_deassert_cnt[1] .is_wysiwyg = "true";
defparam \cs_deassert_cnt[1] .power_up = "low";

cycloneive_lcell_comb \Add5~0 (
	.dataa(\cs_deassert_cnt[0]~q ),
	.datab(\cs_deassert_cnt[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add5~0_combout ),
	.cout());
defparam \Add5~0 .lut_mask = 16'h8888;
defparam \Add5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cs_deassert_cnt_next~5 (
	.dataa(\cs_deassert_cnt[3]~q ),
	.datab(\cs_deassert_cnt[2]~q ),
	.datac(\Add5~0_combout ),
	.datad(\Equal15~3_combout ),
	.cin(gnd),
	.combout(\cs_deassert_cnt_next~5_combout ),
	.cout());
defparam \cs_deassert_cnt_next~5 .lut_mask = 16'h006A;
defparam \cs_deassert_cnt_next~5 .sum_lutc_input = "datac";

dffeas \cs_deassert_cnt[3] (
	.clk(clk_clk),
	.d(\cs_deassert_cnt_next~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.ST_DEASSERT_CS_DLY~q ),
	.q(\cs_deassert_cnt[3]~q ),
	.prn(vcc));
defparam \cs_deassert_cnt[3] .is_wysiwyg = "true";
defparam \cs_deassert_cnt[3] .power_up = "low";

cycloneive_lcell_comb \Equal15~1 (
	.dataa(csr_delay_setting_data_6),
	.datab(\cs_deassert_cnt[2]~q ),
	.datac(csr_delay_setting_data_5),
	.datad(\cs_deassert_cnt[1]~q ),
	.cin(gnd),
	.combout(\Equal15~1_combout ),
	.cout());
defparam \Equal15~1 .lut_mask = 16'h6D66;
defparam \Equal15~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal15~2 (
	.dataa(\cs_deassert_cnt[0]~q ),
	.datab(csr_delay_setting_data_7),
	.datac(\cs_deassert_cnt[3]~q ),
	.datad(\Equal15~1_combout ),
	.cin(gnd),
	.combout(\Equal15~2_combout ),
	.cout());
defparam \Equal15~2 .lut_mask = 16'hD73C;
defparam \Equal15~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cs_deassert_cnt_next~7 (
	.dataa(csr_delay_setting_data_4),
	.datab(\Equal15~0_combout ),
	.datac(\cs_deassert_cnt[0]~q ),
	.datad(\Equal15~2_combout ),
	.cin(gnd),
	.combout(\cs_deassert_cnt_next~7_combout ),
	.cout());
defparam \cs_deassert_cnt_next~7 .lut_mask = 16'h0F0D;
defparam \cs_deassert_cnt_next~7 .sum_lutc_input = "datac";

dffeas \cs_deassert_cnt[0] (
	.clk(clk_clk),
	.d(\cs_deassert_cnt_next~7_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.ST_DEASSERT_CS_DLY~q ),
	.q(\cs_deassert_cnt[0]~q ),
	.prn(vcc));
defparam \cs_deassert_cnt[0] .is_wysiwyg = "true";
defparam \cs_deassert_cnt[0] .power_up = "low";

cycloneive_lcell_comb \cs_deassert_cnt_next~6 (
	.dataa(\cs_deassert_cnt[0]~q ),
	.datab(\cs_deassert_cnt[1]~q ),
	.datac(\cs_deassert_cnt[2]~q ),
	.datad(\Equal15~3_combout ),
	.cin(gnd),
	.combout(\cs_deassert_cnt_next~6_combout ),
	.cout());
defparam \cs_deassert_cnt_next~6 .lut_mask = 16'h0078;
defparam \cs_deassert_cnt_next~6 .sum_lutc_input = "datac";

dffeas \cs_deassert_cnt[2] (
	.clk(clk_clk),
	.d(\cs_deassert_cnt_next~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.ST_DEASSERT_CS_DLY~q ),
	.q(\cs_deassert_cnt[2]~q ),
	.prn(vcc));
defparam \cs_deassert_cnt[2] .is_wysiwyg = "true";
defparam \cs_deassert_cnt[2] .power_up = "low";

cycloneive_lcell_comb \Equal15~0 (
	.dataa(csr_delay_setting_data_6),
	.datab(\cs_deassert_cnt[2]~q ),
	.datac(csr_delay_setting_data_5),
	.datad(\cs_deassert_cnt[1]~q ),
	.cin(gnd),
	.combout(\Equal15~0_combout ),
	.cout());
defparam \Equal15~0 .lut_mask = 16'h0690;
defparam \Equal15~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal15~3 (
	.dataa(csr_delay_setting_data_4),
	.datab(\Equal15~0_combout ),
	.datac(\cs_deassert_cnt[0]~q ),
	.datad(\Equal15~2_combout ),
	.cin(gnd),
	.combout(\Equal15~3_combout ),
	.cout());
defparam \Equal15~3 .lut_mask = 16'h0042;
defparam \Equal15~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector7~0 (
	.dataa(csr_delay_setting_data_4),
	.datab(csr_delay_setting_data_5),
	.datac(csr_delay_setting_data_6),
	.datad(csr_delay_setting_data_7),
	.cin(gnd),
	.combout(\Selector7~0_combout ),
	.cout());
defparam \Selector7~0 .lut_mask = 16'h0001;
defparam \Selector7~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector8~0 (
	.dataa(\state.ST_DEASSERT_CS_DLY~q ),
	.datab(\state.ST_STOP_CLK~q ),
	.datac(\Equal15~3_combout ),
	.datad(\Selector7~0_combout ),
	.cin(gnd),
	.combout(\Selector8~0_combout ),
	.cout());
defparam \Selector8~0 .lut_mask = 16'h0ACE;
defparam \Selector8~0 .sum_lutc_input = "datac";

dffeas \state.ST_DEASSERT_CS_DLY (
	.clk(clk_clk),
	.d(\Selector8~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_DEASSERT_CS_DLY~q ),
	.prn(vcc));
defparam \state.ST_DEASSERT_CS_DLY .is_wysiwyg = "true";
defparam \state.ST_DEASSERT_CS_DLY .power_up = "low";

cycloneive_lcell_comb \Selector7~1 (
	.dataa(\state.ST_DEASSERT_CS_DLY~q ),
	.datab(\state.ST_STOP_CLK~q ),
	.datac(\Selector7~0_combout ),
	.datad(\Equal15~3_combout ),
	.cin(gnd),
	.combout(\Selector7~1_combout ),
	.cout());
defparam \Selector7~1 .lut_mask = 16'hEAC0;
defparam \Selector7~1 .sum_lutc_input = "datac";

dffeas \state.ST_DEASSERT_CS (
	.clk(clk_clk),
	.d(\Selector7~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_DEASSERT_CS~q ),
	.prn(vcc));
defparam \state.ST_DEASSERT_CS .is_wysiwyg = "true";
defparam \state.ST_DEASSERT_CS .power_up = "low";

cycloneive_lcell_comb \ncs_wire[0]~0 (
	.dataa(header_information_30),
	.datab(\state.ST_DEASSERT_CS~q ),
	.datac(\state.ST_IDLE~q ),
	.datad(\state.ST_START_CLK~q ),
	.cin(gnd),
	.combout(\ncs_wire[0]~0_combout ),
	.cout());
defparam \ncs_wire[0]~0 .lut_mask = 16'hAAEF;
defparam \ncs_wire[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ncs_wire[0]~1 (
	.dataa(\ncs_wire[0]~0_combout ),
	.datab(header_information_29),
	.datac(header_information_28),
	.datad(header_information_27),
	.cin(gnd),
	.combout(\ncs_wire[0]~1_combout ),
	.cout());
defparam \ncs_wire[0]~1 .lut_mask = 16'hFFFE;
defparam \ncs_wire[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \ncs_wire[0]~3 (
	.dataa(\ncs_wire[0]~1_combout ),
	.datab(\state.ST_START_CLK~q ),
	.datac(\ncs_wire[0]~2_combout ),
	.datad(csr_delay_setting_data_0),
	.cin(gnd),
	.combout(\ncs_wire[0]~3_combout ),
	.cout());
defparam \ncs_wire[0]~3 .lut_mask = 16'h5515;
defparam \ncs_wire[0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \flash_data_out[0]~0 (
	.dataa(\inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|out_payload[12]~q ),
	.datab(\inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|out_payload[2]~q ),
	.datac(\inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|out_payload[1]~q ),
	.datad(\inf_sc_fifo_ser_data_inst|inf_sc_fifo_ser_data|out_payload[0]~q ),
	.cin(gnd),
	.combout(\flash_data_out[0]~0_combout ),
	.cout());
defparam \flash_data_out[0]~0 .lut_mask = 16'hFEEB;
defparam \flash_data_out[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \demux_channel[2]~0 (
	.dataa(addr_num_lines_2),
	.datab(data_num_lines_2),
	.datac(gnd),
	.datad(stateST_SEND_ADDR),
	.cin(gnd),
	.combout(\demux_channel[2]~0_combout ),
	.cout());
defparam \demux_channel[2]~0 .lut_mask = 16'hAACC;
defparam \demux_channel[2]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(in_cmd_channel_reg_1),
	.datab(gnd),
	.datac(gnd),
	.datad(in_cmd_channel_reg_0),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h00AA;
defparam \Equal0~0 .sum_lutc_input = "datac";

dffeas \read_capture_delay_reg[0] (
	.clk(clk_clk),
	.d(\clk_div_new_inst_2|rising_edge~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(!\state.ST_RECEIVE~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\read_capture_delay_reg[0]~q ),
	.prn(vcc));
defparam \read_capture_delay_reg[0] .is_wysiwyg = "true";
defparam \read_capture_delay_reg[0] .power_up = "low";

cycloneive_lcell_comb \read_capture_delay_reg~9 (
	.dataa(\state.ST_RECEIVE~q ),
	.datab(\read_capture_delay_reg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_capture_delay_reg~9_combout ),
	.cout());
defparam \read_capture_delay_reg~9 .lut_mask = 16'h8888;
defparam \read_capture_delay_reg~9 .sum_lutc_input = "datac";

dffeas \read_capture_delay_reg[1] (
	.clk(clk_clk),
	.d(\read_capture_delay_reg~9_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read_capture_delay_reg[1]~q ),
	.prn(vcc));
defparam \read_capture_delay_reg[1] .is_wysiwyg = "true";
defparam \read_capture_delay_reg[1] .power_up = "low";

cycloneive_lcell_comb \read_capture_delay_reg~8 (
	.dataa(\state.ST_RECEIVE~q ),
	.datab(\read_capture_delay_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_capture_delay_reg~8_combout ),
	.cout());
defparam \read_capture_delay_reg~8 .lut_mask = 16'h8888;
defparam \read_capture_delay_reg~8 .sum_lutc_input = "datac";

dffeas \read_capture_delay_reg[2] (
	.clk(clk_clk),
	.d(\read_capture_delay_reg~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read_capture_delay_reg[2]~q ),
	.prn(vcc));
defparam \read_capture_delay_reg[2] .is_wysiwyg = "true";
defparam \read_capture_delay_reg[2] .power_up = "low";

cycloneive_lcell_comb \read_capture_delay_reg~10 (
	.dataa(\state.ST_RECEIVE~q ),
	.datab(\read_capture_delay_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_capture_delay_reg~10_combout ),
	.cout());
defparam \read_capture_delay_reg~10 .lut_mask = 16'h8888;
defparam \read_capture_delay_reg~10 .sum_lutc_input = "datac";

dffeas \read_capture_delay_reg[3] (
	.clk(clk_clk),
	.d(\read_capture_delay_reg~10_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read_capture_delay_reg[3]~q ),
	.prn(vcc));
defparam \read_capture_delay_reg[3] .is_wysiwyg = "true";
defparam \read_capture_delay_reg[3] .power_up = "low";

cycloneive_lcell_comb \read_capture_delay_reg~6 (
	.dataa(\state.ST_RECEIVE~q ),
	.datab(\read_capture_delay_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_capture_delay_reg~6_combout ),
	.cout());
defparam \read_capture_delay_reg~6 .lut_mask = 16'h8888;
defparam \read_capture_delay_reg~6 .sum_lutc_input = "datac";

dffeas \read_capture_delay_reg[4] (
	.clk(clk_clk),
	.d(\read_capture_delay_reg~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read_capture_delay_reg[4]~q ),
	.prn(vcc));
defparam \read_capture_delay_reg[4] .is_wysiwyg = "true";
defparam \read_capture_delay_reg[4] .power_up = "low";

cycloneive_lcell_comb \read_capture_delay_reg~4 (
	.dataa(\state.ST_RECEIVE~q ),
	.datab(\read_capture_delay_reg[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_capture_delay_reg~4_combout ),
	.cout());
defparam \read_capture_delay_reg~4 .lut_mask = 16'h8888;
defparam \read_capture_delay_reg~4 .sum_lutc_input = "datac";

dffeas \read_capture_delay_reg[5] (
	.clk(clk_clk),
	.d(\read_capture_delay_reg~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read_capture_delay_reg[5]~q ),
	.prn(vcc));
defparam \read_capture_delay_reg[5] .is_wysiwyg = "true";
defparam \read_capture_delay_reg[5] .power_up = "low";

cycloneive_lcell_comb \read_capture_delay_reg~5 (
	.dataa(\state.ST_RECEIVE~q ),
	.datab(\read_capture_delay_reg[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_capture_delay_reg~5_combout ),
	.cout());
defparam \read_capture_delay_reg~5 .lut_mask = 16'h8888;
defparam \read_capture_delay_reg~5 .sum_lutc_input = "datac";

dffeas \read_capture_delay_reg[6] (
	.clk(clk_clk),
	.d(\read_capture_delay_reg~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read_capture_delay_reg[6]~q ),
	.prn(vcc));
defparam \read_capture_delay_reg[6] .is_wysiwyg = "true";
defparam \read_capture_delay_reg[6] .power_up = "low";

cycloneive_lcell_comb \read_capture_delay_reg~7 (
	.dataa(\state.ST_RECEIVE~q ),
	.datab(\read_capture_delay_reg[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_capture_delay_reg~7_combout ),
	.cout());
defparam \read_capture_delay_reg~7 .lut_mask = 16'h8888;
defparam \read_capture_delay_reg~7 .sum_lutc_input = "datac";

dffeas \read_capture_delay_reg[7] (
	.clk(clk_clk),
	.d(\read_capture_delay_reg~7_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read_capture_delay_reg[7]~q ),
	.prn(vcc));
defparam \read_capture_delay_reg[7] .is_wysiwyg = "true";
defparam \read_capture_delay_reg[7] .power_up = "low";

cycloneive_lcell_comb \read_capture_delay_reg~2 (
	.dataa(\state.ST_RECEIVE~q ),
	.datab(\read_capture_delay_reg[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_capture_delay_reg~2_combout ),
	.cout());
defparam \read_capture_delay_reg~2 .lut_mask = 16'h8888;
defparam \read_capture_delay_reg~2 .sum_lutc_input = "datac";

dffeas \read_capture_delay_reg[8] (
	.clk(clk_clk),
	.d(\read_capture_delay_reg~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read_capture_delay_reg[8]~q ),
	.prn(vcc));
defparam \read_capture_delay_reg[8] .is_wysiwyg = "true";
defparam \read_capture_delay_reg[8] .power_up = "low";

cycloneive_lcell_comb \read_capture_delay_reg~1 (
	.dataa(\state.ST_RECEIVE~q ),
	.datab(\read_capture_delay_reg[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_capture_delay_reg~1_combout ),
	.cout());
defparam \read_capture_delay_reg~1 .lut_mask = 16'h8888;
defparam \read_capture_delay_reg~1 .sum_lutc_input = "datac";

dffeas \read_capture_delay_reg[9] (
	.clk(clk_clk),
	.d(\read_capture_delay_reg~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read_capture_delay_reg[9]~q ),
	.prn(vcc));
defparam \read_capture_delay_reg[9] .is_wysiwyg = "true";
defparam \read_capture_delay_reg[9] .power_up = "low";

cycloneive_lcell_comb \read_capture_delay_reg~0 (
	.dataa(\state.ST_RECEIVE~q ),
	.datab(\read_capture_delay_reg[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_capture_delay_reg~0_combout ),
	.cout());
defparam \read_capture_delay_reg~0 .lut_mask = 16'h8888;
defparam \read_capture_delay_reg~0 .sum_lutc_input = "datac";

dffeas \read_capture_delay_reg[10] (
	.clk(clk_clk),
	.d(\read_capture_delay_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read_capture_delay_reg[10]~q ),
	.prn(vcc));
defparam \read_capture_delay_reg[10] .is_wysiwyg = "true";
defparam \read_capture_delay_reg[10] .power_up = "low";

cycloneive_lcell_comb \Mux0~0 (
	.dataa(csr_rd_capturing_data_1),
	.datab(\read_capture_delay_reg[9]~q ),
	.datac(csr_rd_capturing_data_0),
	.datad(\read_capture_delay_reg[8]~q ),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hE5E0;
defparam \Mux0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_capture_delay_reg~3 (
	.dataa(\state.ST_RECEIVE~q ),
	.datab(\read_capture_delay_reg[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_capture_delay_reg~3_combout ),
	.cout());
defparam \read_capture_delay_reg~3 .lut_mask = 16'h8888;
defparam \read_capture_delay_reg~3 .sum_lutc_input = "datac";

dffeas \read_capture_delay_reg[11] (
	.clk(clk_clk),
	.d(\read_capture_delay_reg~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read_capture_delay_reg[11]~q ),
	.prn(vcc));
defparam \read_capture_delay_reg[11] .is_wysiwyg = "true";
defparam \read_capture_delay_reg[11] .power_up = "low";

cycloneive_lcell_comb \Mux0~1 (
	.dataa(\read_capture_delay_reg[10]~q ),
	.datab(csr_rd_capturing_data_1),
	.datac(\Mux0~0_combout ),
	.datad(\read_capture_delay_reg[11]~q ),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hF838;
defparam \Mux0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~2 (
	.dataa(csr_rd_capturing_data_0),
	.datab(\read_capture_delay_reg[6]~q ),
	.datac(csr_rd_capturing_data_1),
	.datad(\read_capture_delay_reg[4]~q ),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
defparam \Mux0~2 .lut_mask = 16'hE5E0;
defparam \Mux0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~3 (
	.dataa(\read_capture_delay_reg[5]~q ),
	.datab(csr_rd_capturing_data_0),
	.datac(\Mux0~2_combout ),
	.datad(\read_capture_delay_reg[7]~q ),
	.cin(gnd),
	.combout(\Mux0~3_combout ),
	.cout());
defparam \Mux0~3 .lut_mask = 16'hF838;
defparam \Mux0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~4 (
	.dataa(csr_rd_capturing_data_1),
	.datab(\read_capture_delay_reg[1]~q ),
	.datac(csr_rd_capturing_data_0),
	.datad(\read_capture_delay_reg[0]~q ),
	.cin(gnd),
	.combout(\Mux0~4_combout ),
	.cout());
defparam \Mux0~4 .lut_mask = 16'hE5E0;
defparam \Mux0~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~5 (
	.dataa(\read_capture_delay_reg[2]~q ),
	.datab(csr_rd_capturing_data_1),
	.datac(\Mux0~4_combout ),
	.datad(\read_capture_delay_reg[3]~q ),
	.cin(gnd),
	.combout(\Mux0~5_combout ),
	.cout());
defparam \Mux0~5 .lut_mask = 16'hF838;
defparam \Mux0~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~6 (
	.dataa(csr_rd_capturing_data_3),
	.datab(\Mux0~3_combout ),
	.datac(csr_rd_capturing_data_2),
	.datad(\Mux0~5_combout ),
	.cin(gnd),
	.combout(\Mux0~6_combout ),
	.cout());
defparam \Mux0~6 .lut_mask = 16'hE5E0;
defparam \Mux0~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_capture_delay_reg~12 (
	.dataa(\state.ST_RECEIVE~q ),
	.datab(\read_capture_delay_reg[11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_capture_delay_reg~12_combout ),
	.cout());
defparam \read_capture_delay_reg~12 .lut_mask = 16'h8888;
defparam \read_capture_delay_reg~12 .sum_lutc_input = "datac";

dffeas \read_capture_delay_reg[12] (
	.clk(clk_clk),
	.d(\read_capture_delay_reg~12_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read_capture_delay_reg[12]~q ),
	.prn(vcc));
defparam \read_capture_delay_reg[12] .is_wysiwyg = "true";
defparam \read_capture_delay_reg[12] .power_up = "low";

cycloneive_lcell_comb \read_capture_delay_reg~11 (
	.dataa(\state.ST_RECEIVE~q ),
	.datab(\read_capture_delay_reg[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_capture_delay_reg~11_combout ),
	.cout());
defparam \read_capture_delay_reg~11 .lut_mask = 16'h8888;
defparam \read_capture_delay_reg~11 .sum_lutc_input = "datac";

dffeas \read_capture_delay_reg[13] (
	.clk(clk_clk),
	.d(\read_capture_delay_reg~11_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read_capture_delay_reg[13]~q ),
	.prn(vcc));
defparam \read_capture_delay_reg[13] .is_wysiwyg = "true";
defparam \read_capture_delay_reg[13] .power_up = "low";

cycloneive_lcell_comb \Mux0~7 (
	.dataa(\read_capture_delay_reg[13]~q ),
	.datab(\read_capture_delay_reg[12]~q ),
	.datac(csr_rd_capturing_data_0),
	.datad(csr_rd_capturing_data_1),
	.cin(gnd),
	.combout(\Mux0~7_combout ),
	.cout());
defparam \Mux0~7 .lut_mask = 16'h00AC;
defparam \Mux0~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_capture_delay_reg~13 (
	.dataa(\state.ST_RECEIVE~q ),
	.datab(\read_capture_delay_reg[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_capture_delay_reg~13_combout ),
	.cout());
defparam \read_capture_delay_reg~13 .lut_mask = 16'h8888;
defparam \read_capture_delay_reg~13 .sum_lutc_input = "datac";

dffeas \read_capture_delay_reg[14] (
	.clk(clk_clk),
	.d(\read_capture_delay_reg~13_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read_capture_delay_reg[14]~q ),
	.prn(vcc));
defparam \read_capture_delay_reg[14] .is_wysiwyg = "true";
defparam \read_capture_delay_reg[14] .power_up = "low";

cycloneive_lcell_comb \Mux0~8 (
	.dataa(\Mux0~7_combout ),
	.datab(csr_rd_capturing_data_1),
	.datac(\read_capture_delay_reg[14]~q ),
	.datad(csr_rd_capturing_data_0),
	.cin(gnd),
	.combout(\Mux0~8_combout ),
	.cout());
defparam \Mux0~8 .lut_mask = 16'hAAEA;
defparam \Mux0~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~9 (
	.dataa(\Mux0~1_combout ),
	.datab(csr_rd_capturing_data_3),
	.datac(\Mux0~6_combout ),
	.datad(\Mux0~8_combout ),
	.cin(gnd),
	.combout(\Mux0~9_combout ),
	.cout());
defparam \Mux0~9 .lut_mask = 16'hF838;
defparam \Mux0~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal16~0 (
	.dataa(data_num_lines_0),
	.datab(gnd),
	.datac(data_num_lines_2),
	.datad(data_num_lines_1),
	.cin(gnd),
	.combout(\Equal16~0_combout ),
	.cout());
defparam \Equal16~0 .lut_mask = 16'h000A;
defparam \Equal16~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_data_cnt~2 (
	.dataa(gnd),
	.datab(data_num_lines_0),
	.datac(data_num_lines_1),
	.datad(data_num_lines_2),
	.cin(gnd),
	.combout(\read_data_cnt~2_combout ),
	.cout());
defparam \read_data_cnt~2 .lut_mask = 16'h003C;
defparam \read_data_cnt~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_data_cnt~4 (
	.dataa(\state.ST_SEND~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\read_data_cnt[0]~q ),
	.cin(gnd),
	.combout(\read_data_cnt~4_combout ),
	.cout());
defparam \read_data_cnt~4 .lut_mask = 16'hAAFF;
defparam \read_data_cnt~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_data_cnt[0]~1 (
	.dataa(\state.ST_SEND~q ),
	.datab(\state.ST_RECEIVE~q ),
	.datac(\Mux0~9_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_data_cnt[0]~1_combout ),
	.cout());
defparam \read_data_cnt[0]~1 .lut_mask = 16'hEAEA;
defparam \read_data_cnt[0]~1 .sum_lutc_input = "datac";

dffeas \read_data_cnt[0] (
	.clk(clk_clk),
	.d(\read_data_cnt~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_cnt[0]~1_combout ),
	.q(\read_data_cnt[0]~q ),
	.prn(vcc));
defparam \read_data_cnt[0] .is_wysiwyg = "true";
defparam \read_data_cnt[0] .power_up = "low";

cycloneive_lcell_comb \Add6~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\read_data_cnt[1]~q ),
	.datad(\read_data_cnt[0]~q ),
	.cin(gnd),
	.combout(\Add6~1_combout ),
	.cout());
defparam \Add6~1 .lut_mask = 16'h0FF0;
defparam \Add6~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_data_cnt~3 (
	.dataa(\read_data_cnt~2_combout ),
	.datab(\state.ST_SEND~q ),
	.datac(\read_data_done~combout ),
	.datad(\Add6~1_combout ),
	.cin(gnd),
	.combout(\read_data_cnt~3_combout ),
	.cout());
defparam \read_data_cnt~3 .lut_mask = 16'hA8AB;
defparam \read_data_cnt~3 .sum_lutc_input = "datac";

dffeas \read_data_cnt[1] (
	.clk(clk_clk),
	.d(\read_data_cnt~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_cnt[0]~1_combout ),
	.q(\read_data_cnt[1]~q ),
	.prn(vcc));
defparam \read_data_cnt[1] .is_wysiwyg = "true";
defparam \read_data_cnt[1] .power_up = "low";

cycloneive_lcell_comb \Add6~0 (
	.dataa(gnd),
	.datab(\read_data_cnt[1]~q ),
	.datac(\read_data_cnt[0]~q ),
	.datad(\read_data_cnt[2]~q ),
	.cin(gnd),
	.combout(\Add6~0_combout ),
	.cout());
defparam \Add6~0 .lut_mask = 16'h03FC;
defparam \Add6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_data_cnt~0 (
	.dataa(\Equal16~0_combout ),
	.datab(\state.ST_SEND~q ),
	.datac(\read_data_done~combout ),
	.datad(\Add6~0_combout ),
	.cin(gnd),
	.combout(\read_data_cnt~0_combout ),
	.cout());
defparam \read_data_cnt~0 .lut_mask = 16'hA8AB;
defparam \read_data_cnt~0 .sum_lutc_input = "datac";

dffeas \read_data_cnt[2] (
	.clk(clk_clk),
	.d(\read_data_cnt~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_cnt[0]~1_combout ),
	.q(\read_data_cnt[2]~q ),
	.prn(vcc));
defparam \read_data_cnt[2] .is_wysiwyg = "true";
defparam \read_data_cnt[2] .power_up = "low";

cycloneive_lcell_comb \read_data_done~0 (
	.dataa(gnd),
	.datab(\read_data_cnt[2]~q ),
	.datac(\read_data_cnt[1]~q ),
	.datad(\read_data_cnt[0]~q ),
	.cin(gnd),
	.combout(\read_data_done~0_combout ),
	.cout());
defparam \read_data_done~0 .lut_mask = 16'h0003;
defparam \read_data_done~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_data_cnt~5 (
	.dataa(\state.ST_SEND~q ),
	.datab(\read_data_done~combout ),
	.datac(\read_data_cnt[3]~q ),
	.datad(\read_data_done~0_combout ),
	.cin(gnd),
	.combout(\read_data_cnt~5_combout ),
	.cout());
defparam \read_data_cnt~5 .lut_mask = 16'h0110;
defparam \read_data_cnt~5 .sum_lutc_input = "datac";

dffeas \read_data_cnt[3] (
	.clk(clk_clk),
	.d(\read_data_cnt~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_cnt[0]~1_combout ),
	.q(\read_data_cnt[3]~q ),
	.prn(vcc));
defparam \read_data_cnt[3] .is_wysiwyg = "true";
defparam \read_data_cnt[3] .power_up = "low";

cycloneive_lcell_comb read_data_done(
	.dataa(\state.ST_RECEIVE~q ),
	.datab(\Mux0~9_combout ),
	.datac(\read_data_done~0_combout ),
	.datad(\read_data_cnt[3]~q ),
	.cin(gnd),
	.combout(\read_data_done~combout ),
	.cout());
defparam read_data_done.lut_mask = 16'h0080;
defparam read_data_done.sum_lutc_input = "datac";

dffeas read_data_valid(
	.clk(clk_clk),
	.d(\read_data_done~combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read_data_valid~q ),
	.prn(vcc));
defparam read_data_valid.is_wysiwyg = "true";
defparam read_data_valid.power_up = "low";

cycloneive_lcell_comb \flash_datain_reg~4 (
	.dataa(data_num_lines_0),
	.datab(dut_asmiblock),
	.datac(data_num_lines_2),
	.datad(data_num_lines_1),
	.cin(gnd),
	.combout(\flash_datain_reg~4_combout ),
	.cout());
defparam \flash_datain_reg~4 .lut_mask = 16'h0008;
defparam \flash_datain_reg~4 .sum_lutc_input = "datac";

dffeas \flash_datain_reg[0] (
	.clk(clk_clk),
	.d(\flash_datain_reg~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux0~9_combout ),
	.q(\flash_datain_reg[0]~q ),
	.prn(vcc));
defparam \flash_datain_reg[0] .is_wysiwyg = "true";
defparam \flash_datain_reg[0] .power_up = "low";

cycloneive_lcell_comb \flash_datain_reg~5 (
	.dataa(\flash_datain_reg[0]~q ),
	.datab(dut_asmiblock),
	.datac(gnd),
	.datad(\Equal16~0_combout ),
	.cin(gnd),
	.combout(\flash_datain_reg~5_combout ),
	.cout());
defparam \flash_datain_reg~5 .lut_mask = 16'hAACC;
defparam \flash_datain_reg~5 .sum_lutc_input = "datac";

dffeas \flash_datain_reg[1] (
	.clk(clk_clk),
	.d(\flash_datain_reg~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux0~9_combout ),
	.q(\flash_datain_reg[1]~q ),
	.prn(vcc));
defparam \flash_datain_reg[1] .is_wysiwyg = "true";
defparam \flash_datain_reg[1] .power_up = "low";

cycloneive_lcell_comb \Equal17~0 (
	.dataa(data_num_lines_1),
	.datab(gnd),
	.datac(data_num_lines_2),
	.datad(data_num_lines_0),
	.cin(gnd),
	.combout(\Equal17~0_combout ),
	.cout());
defparam \Equal17~0 .lut_mask = 16'h000A;
defparam \Equal17~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \flash_datain_reg~6 (
	.dataa(\flash_datain_reg[1]~q ),
	.datab(\flash_datain_reg[0]~q ),
	.datac(\Equal17~0_combout ),
	.datad(\Equal16~0_combout ),
	.cin(gnd),
	.combout(\flash_datain_reg~6_combout ),
	.cout());
defparam \flash_datain_reg~6 .lut_mask = 16'hAAC0;
defparam \flash_datain_reg~6 .sum_lutc_input = "datac";

dffeas \flash_datain_reg[2] (
	.clk(clk_clk),
	.d(\flash_datain_reg~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux0~9_combout ),
	.q(\flash_datain_reg[2]~q ),
	.prn(vcc));
defparam \flash_datain_reg[2] .is_wysiwyg = "true";
defparam \flash_datain_reg[2] .power_up = "low";

cycloneive_lcell_comb \flash_datain_reg~7 (
	.dataa(\flash_datain_reg[2]~q ),
	.datab(\flash_datain_reg[1]~q ),
	.datac(\Equal17~0_combout ),
	.datad(\Equal16~0_combout ),
	.cin(gnd),
	.combout(\flash_datain_reg~7_combout ),
	.cout());
defparam \flash_datain_reg~7 .lut_mask = 16'hAAC0;
defparam \flash_datain_reg~7 .sum_lutc_input = "datac";

dffeas \flash_datain_reg[3] (
	.clk(clk_clk),
	.d(\flash_datain_reg~7_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Mux0~9_combout ),
	.q(\flash_datain_reg[3]~q ),
	.prn(vcc));
defparam \flash_datain_reg[3] .is_wysiwyg = "true";
defparam \flash_datain_reg[3] .power_up = "low";

cycloneive_lcell_comb \flash_datain_reg[4]~0 (
	.dataa(\flash_datain_reg[0]~q ),
	.datab(\flash_datain_reg[2]~q ),
	.datac(gnd),
	.datad(\Equal17~0_combout ),
	.cin(gnd),
	.combout(\flash_datain_reg[4]~0_combout ),
	.cout());
defparam \flash_datain_reg[4]~0 .lut_mask = 16'hCCAA;
defparam \flash_datain_reg[4]~0 .sum_lutc_input = "datac";

dffeas \flash_datain_reg[4] (
	.clk(clk_clk),
	.d(\flash_datain_reg[4]~0_combout ),
	.asdata(\flash_datain_reg[3]~q ),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal16~0_combout ),
	.ena(\Mux0~9_combout ),
	.q(\flash_datain_reg[4]~q ),
	.prn(vcc));
defparam \flash_datain_reg[4] .is_wysiwyg = "true";
defparam \flash_datain_reg[4] .power_up = "low";

cycloneive_lcell_comb \flash_datain_reg[5]~1 (
	.dataa(\flash_datain_reg[1]~q ),
	.datab(\flash_datain_reg[3]~q ),
	.datac(gnd),
	.datad(\Equal17~0_combout ),
	.cin(gnd),
	.combout(\flash_datain_reg[5]~1_combout ),
	.cout());
defparam \flash_datain_reg[5]~1 .lut_mask = 16'hCCAA;
defparam \flash_datain_reg[5]~1 .sum_lutc_input = "datac";

dffeas \flash_datain_reg[5] (
	.clk(clk_clk),
	.d(\flash_datain_reg[5]~1_combout ),
	.asdata(\flash_datain_reg[4]~q ),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal16~0_combout ),
	.ena(\Mux0~9_combout ),
	.q(\flash_datain_reg[5]~q ),
	.prn(vcc));
defparam \flash_datain_reg[5] .is_wysiwyg = "true";
defparam \flash_datain_reg[5] .power_up = "low";

cycloneive_lcell_comb \flash_datain_reg[6]~2 (
	.dataa(\flash_datain_reg[2]~q ),
	.datab(\flash_datain_reg[4]~q ),
	.datac(gnd),
	.datad(\Equal17~0_combout ),
	.cin(gnd),
	.combout(\flash_datain_reg[6]~2_combout ),
	.cout());
defparam \flash_datain_reg[6]~2 .lut_mask = 16'hCCAA;
defparam \flash_datain_reg[6]~2 .sum_lutc_input = "datac";

dffeas \flash_datain_reg[6] (
	.clk(clk_clk),
	.d(\flash_datain_reg[6]~2_combout ),
	.asdata(\flash_datain_reg[5]~q ),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal16~0_combout ),
	.ena(\Mux0~9_combout ),
	.q(\flash_datain_reg[6]~q ),
	.prn(vcc));
defparam \flash_datain_reg[6] .is_wysiwyg = "true";
defparam \flash_datain_reg[6] .power_up = "low";

cycloneive_lcell_comb \flash_datain_reg[7]~3 (
	.dataa(\flash_datain_reg[3]~q ),
	.datab(\flash_datain_reg[5]~q ),
	.datac(gnd),
	.datad(\Equal17~0_combout ),
	.cin(gnd),
	.combout(\flash_datain_reg[7]~3_combout ),
	.cout());
defparam \flash_datain_reg[7]~3 .lut_mask = 16'hCCAA;
defparam \flash_datain_reg[7]~3 .sum_lutc_input = "datac";

dffeas \flash_datain_reg[7] (
	.clk(clk_clk),
	.d(\flash_datain_reg[7]~3_combout ),
	.asdata(\flash_datain_reg[6]~q ),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal16~0_combout ),
	.ena(\Mux0~9_combout ),
	.q(\flash_datain_reg[7]~q ),
	.prn(vcc));
defparam \flash_datain_reg[7] .is_wysiwyg = "true";
defparam \flash_datain_reg[7] .power_up = "low";

endmodule

module flashLoader_adapter_8_1 (
	reset_n,
	in_channel,
	grant_0,
	out_valid1,
	full_addercout_1,
	cout,
	mem_used_9,
	in_ready1,
	grant_01,
	out_endofpacket1,
	in_valid,
	out_data_0,
	out_channel_2,
	out_channel_1,
	out_channel_0,
	out_channel_8,
	in_endofpacket,
	in_data,
	clk)/* synthesis synthesis_greybox=0 */;
input 	reset_n;
input 	[11:0] in_channel;
input 	grant_0;
output 	out_valid1;
input 	full_addercout_1;
input 	cout;
input 	mem_used_9;
output 	in_ready1;
input 	grant_01;
output 	out_endofpacket1;
input 	in_valid;
output 	out_data_0;
output 	out_channel_2;
output 	out_channel_1;
output 	out_channel_0;
output 	out_channel_8;
input 	in_endofpacket;
input 	[7:0] in_data;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a_valid~q ;
wire \always4~1_combout ;
wire \always4~0_combout ;
wire \state_register[0]~0_combout ;
wire \state_register[0]~q ;
wire \Mux3~0_combout ;
wire \state_register[1]~q ;
wire \Mux2~0_combout ;
wire \Mux2~1_combout ;
wire \state_register[2]~q ;
wire \Mux1~0_combout ;
wire \a_endofpacket~q ;
wire \Mux5~0_combout ;
wire \a_data5[0]~q ;
wire \a_data6[0]~q ;
wire \a_data4[0]~q ;
wire \Mux0~0_combout ;
wire \a_data7[0]~q ;
wire \Mux0~1_combout ;
wire \a_data2[0]~q ;
wire \a_data1[0]~q ;
wire \a_data0[0]~q ;
wire \Mux0~2_combout ;
wire \a_data3[0]~q ;
wire \Mux0~3_combout ;
wire \Mux0~4_combout ;
wire \a_channel[2]~q ;
wire \a_channel[1]~q ;
wire \a_channel[0]~q ;
wire \a_channel[8]~q ;


dffeas out_valid(
	.clk(clk),
	.d(\a_valid~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~1_combout ),
	.q(out_valid1),
	.prn(vcc));
defparam out_valid.is_wysiwyg = "true";
defparam out_valid.power_up = "low";

cycloneive_lcell_comb in_ready(
	.dataa(\Mux1~0_combout ),
	.datab(\always4~0_combout ),
	.datac(out_valid1),
	.datad(\a_valid~q ),
	.cin(gnd),
	.combout(in_ready1),
	.cout());
defparam in_ready.lut_mask = 16'h8AFF;
defparam in_ready.sum_lutc_input = "datac";

dffeas out_endofpacket(
	.clk(clk),
	.d(\Mux5~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~1_combout ),
	.q(out_endofpacket1),
	.prn(vcc));
defparam out_endofpacket.is_wysiwyg = "true";
defparam out_endofpacket.power_up = "low";

dffeas \out_data[0] (
	.clk(clk),
	.d(\Mux0~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~1_combout ),
	.q(out_data_0),
	.prn(vcc));
defparam \out_data[0] .is_wysiwyg = "true";
defparam \out_data[0] .power_up = "low";

dffeas \out_channel[2] (
	.clk(clk),
	.d(\a_channel[2]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~1_combout ),
	.q(out_channel_2),
	.prn(vcc));
defparam \out_channel[2] .is_wysiwyg = "true";
defparam \out_channel[2] .power_up = "low";

dffeas \out_channel[1] (
	.clk(clk),
	.d(\a_channel[1]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~1_combout ),
	.q(out_channel_1),
	.prn(vcc));
defparam \out_channel[1] .is_wysiwyg = "true";
defparam \out_channel[1] .power_up = "low";

dffeas \out_channel[0] (
	.clk(clk),
	.d(\a_channel[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~1_combout ),
	.q(out_channel_0),
	.prn(vcc));
defparam \out_channel[0] .is_wysiwyg = "true";
defparam \out_channel[0] .power_up = "low";

dffeas \out_channel[8] (
	.clk(clk),
	.d(\a_channel[8]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~1_combout ),
	.q(out_channel_8),
	.prn(vcc));
defparam \out_channel[8] .is_wysiwyg = "true";
defparam \out_channel[8] .power_up = "low";

dffeas a_valid(
	.clk(clk),
	.d(in_valid),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_valid~q ),
	.prn(vcc));
defparam a_valid.is_wysiwyg = "true";
defparam a_valid.power_up = "low";

cycloneive_lcell_comb \always4~1 (
	.dataa(grant_01),
	.datab(gnd),
	.datac(mem_used_9),
	.datad(out_valid1),
	.cin(gnd),
	.combout(\always4~1_combout ),
	.cout());
defparam \always4~1 .lut_mask = 16'h0AFF;
defparam \always4~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always4~0 (
	.dataa(grant_0),
	.datab(full_addercout_1),
	.datac(cout),
	.datad(mem_used_9),
	.cin(gnd),
	.combout(\always4~0_combout ),
	.cout());
defparam \always4~0 .lut_mask = 16'h00AE;
defparam \always4~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \state_register[0]~0 (
	.dataa(out_valid1),
	.datab(\always4~0_combout ),
	.datac(\state_register[0]~q ),
	.datad(\a_valid~q ),
	.cin(gnd),
	.combout(\state_register[0]~0_combout ),
	.cout());
defparam \state_register[0]~0 .lut_mask = 16'h2DF0;
defparam \state_register[0]~0 .sum_lutc_input = "datac";

dffeas \state_register[0] (
	.clk(clk),
	.d(\state_register[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state_register[0]~q ),
	.prn(vcc));
defparam \state_register[0] .is_wysiwyg = "true";
defparam \state_register[0] .power_up = "low";

cycloneive_lcell_comb \Mux3~0 (
	.dataa(\state_register[1]~q ),
	.datab(\a_valid~q ),
	.datac(\always4~1_combout ),
	.datad(\state_register[0]~q ),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'h6AAA;
defparam \Mux3~0 .sum_lutc_input = "datac";

dffeas \state_register[1] (
	.clk(clk),
	.d(\Mux3~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state_register[1]~q ),
	.prn(vcc));
defparam \state_register[1] .is_wysiwyg = "true";
defparam \state_register[1] .power_up = "low";

cycloneive_lcell_comb \Mux2~0 (
	.dataa(\a_valid~q ),
	.datab(\state_register[0]~q ),
	.datac(\always4~0_combout ),
	.datad(out_valid1),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
defparam \Mux2~0 .lut_mask = 16'h8088;
defparam \Mux2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux2~1 (
	.dataa(gnd),
	.datab(\state_register[2]~q ),
	.datac(\state_register[1]~q ),
	.datad(\Mux2~0_combout ),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
defparam \Mux2~1 .lut_mask = 16'h3CCC;
defparam \Mux2~1 .sum_lutc_input = "datac";

dffeas \state_register[2] (
	.clk(clk),
	.d(\Mux2~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state_register[2]~q ),
	.prn(vcc));
defparam \state_register[2] .is_wysiwyg = "true";
defparam \state_register[2] .power_up = "low";

cycloneive_lcell_comb \Mux1~0 (
	.dataa(\state_register[2]~q ),
	.datab(\state_register[1]~q ),
	.datac(\state_register[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'h8080;
defparam \Mux1~0 .sum_lutc_input = "datac";

dffeas a_endofpacket(
	.clk(clk),
	.d(in_endofpacket),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_endofpacket~q ),
	.prn(vcc));
defparam a_endofpacket.is_wysiwyg = "true";
defparam a_endofpacket.power_up = "low";

cycloneive_lcell_comb \Mux5~0 (
	.dataa(\a_valid~q ),
	.datab(\Mux1~0_combout ),
	.datac(\a_endofpacket~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
defparam \Mux5~0 .lut_mask = 16'h8080;
defparam \Mux5~0 .sum_lutc_input = "datac";

dffeas \a_data5[0] (
	.clk(clk),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_data5[0]~q ),
	.prn(vcc));
defparam \a_data5[0] .is_wysiwyg = "true";
defparam \a_data5[0] .power_up = "low";

dffeas \a_data6[0] (
	.clk(clk),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_data6[0]~q ),
	.prn(vcc));
defparam \a_data6[0] .is_wysiwyg = "true";
defparam \a_data6[0] .power_up = "low";

dffeas \a_data4[0] (
	.clk(clk),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_data4[0]~q ),
	.prn(vcc));
defparam \a_data4[0] .is_wysiwyg = "true";
defparam \a_data4[0] .power_up = "low";

cycloneive_lcell_comb \Mux0~0 (
	.dataa(\state_register[0]~q ),
	.datab(\a_data6[0]~q ),
	.datac(\state_register[1]~q ),
	.datad(\a_data4[0]~q ),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hE5E0;
defparam \Mux0~0 .sum_lutc_input = "datac";

dffeas \a_data7[0] (
	.clk(clk),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_data7[0]~q ),
	.prn(vcc));
defparam \a_data7[0] .is_wysiwyg = "true";
defparam \a_data7[0] .power_up = "low";

cycloneive_lcell_comb \Mux0~1 (
	.dataa(\a_data5[0]~q ),
	.datab(\state_register[0]~q ),
	.datac(\Mux0~0_combout ),
	.datad(\a_data7[0]~q ),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hF838;
defparam \Mux0~1 .sum_lutc_input = "datac";

dffeas \a_data2[0] (
	.clk(clk),
	.d(in_data[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_data2[0]~q ),
	.prn(vcc));
defparam \a_data2[0] .is_wysiwyg = "true";
defparam \a_data2[0] .power_up = "low";

dffeas \a_data1[0] (
	.clk(clk),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_data1[0]~q ),
	.prn(vcc));
defparam \a_data1[0] .is_wysiwyg = "true";
defparam \a_data1[0] .power_up = "low";

dffeas \a_data0[0] (
	.clk(clk),
	.d(in_data[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_data0[0]~q ),
	.prn(vcc));
defparam \a_data0[0] .is_wysiwyg = "true";
defparam \a_data0[0] .power_up = "low";

cycloneive_lcell_comb \Mux0~2 (
	.dataa(\state_register[1]~q ),
	.datab(\a_data1[0]~q ),
	.datac(\state_register[0]~q ),
	.datad(\a_data0[0]~q ),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
defparam \Mux0~2 .lut_mask = 16'hE5E0;
defparam \Mux0~2 .sum_lutc_input = "datac";

dffeas \a_data3[0] (
	.clk(clk),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_data3[0]~q ),
	.prn(vcc));
defparam \a_data3[0] .is_wysiwyg = "true";
defparam \a_data3[0] .power_up = "low";

cycloneive_lcell_comb \Mux0~3 (
	.dataa(\a_data2[0]~q ),
	.datab(\state_register[1]~q ),
	.datac(\Mux0~2_combout ),
	.datad(\a_data3[0]~q ),
	.cin(gnd),
	.combout(\Mux0~3_combout ),
	.cout());
defparam \Mux0~3 .lut_mask = 16'hF838;
defparam \Mux0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux0~4 (
	.dataa(\Mux0~1_combout ),
	.datab(\Mux0~3_combout ),
	.datac(gnd),
	.datad(\state_register[2]~q ),
	.cin(gnd),
	.combout(\Mux0~4_combout ),
	.cout());
defparam \Mux0~4 .lut_mask = 16'hAACC;
defparam \Mux0~4 .sum_lutc_input = "datac";

dffeas \a_channel[2] (
	.clk(clk),
	.d(in_channel[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_channel[2]~q ),
	.prn(vcc));
defparam \a_channel[2] .is_wysiwyg = "true";
defparam \a_channel[2] .power_up = "low";

dffeas \a_channel[1] (
	.clk(clk),
	.d(in_channel[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_channel[1]~q ),
	.prn(vcc));
defparam \a_channel[1] .is_wysiwyg = "true";
defparam \a_channel[1] .power_up = "low";

dffeas \a_channel[0] (
	.clk(clk),
	.d(in_channel[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_channel[0]~q ),
	.prn(vcc));
defparam \a_channel[0] .is_wysiwyg = "true";
defparam \a_channel[0] .power_up = "low";

dffeas \a_channel[8] (
	.clk(clk),
	.d(in_channel[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_channel[8]~q ),
	.prn(vcc));
defparam \a_channel[8] .is_wysiwyg = "true";
defparam \a_channel[8] .power_up = "low";

endmodule

module flashLoader_adapter_8_2 (
	reset_n,
	in_channel,
	out_valid1,
	request_1,
	mem_used_9,
	state_register_1,
	state_register_0,
	a_valid1,
	sum_1,
	cout,
	always4,
	in_ready1,
	out_endofpacket1,
	in_valid,
	out_data_0,
	out_channel_2,
	out_channel_1,
	out_channel_0,
	out_channel_8,
	in_endofpacket,
	in_data,
	clk)/* synthesis synthesis_greybox=0 */;
input 	reset_n;
input 	[11:0] in_channel;
output 	out_valid1;
input 	request_1;
input 	mem_used_9;
output 	state_register_1;
output 	state_register_0;
output 	a_valid1;
input 	sum_1;
input 	cout;
output 	always4;
output 	in_ready1;
output 	out_endofpacket1;
input 	in_valid;
output 	out_data_0;
output 	out_channel_2;
output 	out_channel_1;
output 	out_channel_0;
output 	out_channel_8;
input 	in_endofpacket;
input 	[7:0] in_data;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mux4~0_combout ;
wire \state_register[0]~0_combout ;
wire \always4~0_combout ;
wire \a_endofpacket~q ;
wire \Mux6~0_combout ;
wire \a_data5[0]~q ;
wire \a_data3[0]~q ;
wire \a_data1[0]~q ;
wire \Mux1~0_combout ;
wire \a_data7[0]~q ;
wire \Mux1~1_combout ;
wire \a_channel[2]~q ;
wire \a_channel[1]~q ;
wire \a_channel[0]~q ;
wire \a_channel[8]~q ;


dffeas out_valid(
	.clk(clk),
	.d(a_valid1),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always4),
	.q(out_valid1),
	.prn(vcc));
defparam out_valid.is_wysiwyg = "true";
defparam out_valid.power_up = "low";

dffeas \state_register[1] (
	.clk(clk),
	.d(\Mux4~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(state_register_1),
	.prn(vcc));
defparam \state_register[1] .is_wysiwyg = "true";
defparam \state_register[1] .power_up = "low";

dffeas \state_register[0] (
	.clk(clk),
	.d(\state_register[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(state_register_0),
	.prn(vcc));
defparam \state_register[0] .is_wysiwyg = "true";
defparam \state_register[0] .power_up = "low";

dffeas a_valid(
	.clk(clk),
	.d(in_valid),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(a_valid1),
	.prn(vcc));
defparam a_valid.is_wysiwyg = "true";
defparam a_valid.power_up = "low";

cycloneive_lcell_comb \always4~1 (
	.dataa(\always4~0_combout ),
	.datab(request_1),
	.datac(cout),
	.datad(mem_used_9),
	.cin(gnd),
	.combout(always4),
	.cout());
defparam \always4~1 .lut_mask = 16'hAAEB;
defparam \always4~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb in_ready(
	.dataa(state_register_1),
	.datab(state_register_0),
	.datac(always4),
	.datad(a_valid1),
	.cin(gnd),
	.combout(in_ready1),
	.cout());
defparam in_ready.lut_mask = 16'h80FF;
defparam in_ready.sum_lutc_input = "datac";

dffeas out_endofpacket(
	.clk(clk),
	.d(\Mux6~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always4),
	.q(out_endofpacket1),
	.prn(vcc));
defparam out_endofpacket.is_wysiwyg = "true";
defparam out_endofpacket.power_up = "low";

dffeas \out_data[0] (
	.clk(clk),
	.d(\Mux1~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always4),
	.q(out_data_0),
	.prn(vcc));
defparam \out_data[0] .is_wysiwyg = "true";
defparam \out_data[0] .power_up = "low";

dffeas \out_channel[2] (
	.clk(clk),
	.d(\a_channel[2]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always4),
	.q(out_channel_2),
	.prn(vcc));
defparam \out_channel[2] .is_wysiwyg = "true";
defparam \out_channel[2] .power_up = "low";

dffeas \out_channel[1] (
	.clk(clk),
	.d(\a_channel[1]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always4),
	.q(out_channel_1),
	.prn(vcc));
defparam \out_channel[1] .is_wysiwyg = "true";
defparam \out_channel[1] .power_up = "low";

dffeas \out_channel[0] (
	.clk(clk),
	.d(\a_channel[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always4),
	.q(out_channel_0),
	.prn(vcc));
defparam \out_channel[0] .is_wysiwyg = "true";
defparam \out_channel[0] .power_up = "low";

dffeas \out_channel[8] (
	.clk(clk),
	.d(\a_channel[8]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always4),
	.q(out_channel_8),
	.prn(vcc));
defparam \out_channel[8] .is_wysiwyg = "true";
defparam \out_channel[8] .power_up = "low";

cycloneive_lcell_comb \Mux4~0 (
	.dataa(state_register_1),
	.datab(a_valid1),
	.datac(state_register_0),
	.datad(always4),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
defparam \Mux4~0 .lut_mask = 16'h6AAA;
defparam \Mux4~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \state_register[0]~0 (
	.dataa(gnd),
	.datab(state_register_0),
	.datac(a_valid1),
	.datad(always4),
	.cin(gnd),
	.combout(\state_register[0]~0_combout ),
	.cout());
defparam \state_register[0]~0 .lut_mask = 16'h3CCC;
defparam \state_register[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always4~0 (
	.dataa(gnd),
	.datab(mem_used_9),
	.datac(sum_1),
	.datad(out_valid1),
	.cin(gnd),
	.combout(\always4~0_combout ),
	.cout());
defparam \always4~0 .lut_mask = 16'h03FF;
defparam \always4~0 .sum_lutc_input = "datac";

dffeas a_endofpacket(
	.clk(clk),
	.d(in_endofpacket),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_endofpacket~q ),
	.prn(vcc));
defparam a_endofpacket.is_wysiwyg = "true";
defparam a_endofpacket.power_up = "low";

cycloneive_lcell_comb \Mux6~0 (
	.dataa(a_valid1),
	.datab(state_register_1),
	.datac(state_register_0),
	.datad(\a_endofpacket~q ),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
defparam \Mux6~0 .lut_mask = 16'h8000;
defparam \Mux6~0 .sum_lutc_input = "datac";

dffeas \a_data5[0] (
	.clk(clk),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_data5[0]~q ),
	.prn(vcc));
defparam \a_data5[0] .is_wysiwyg = "true";
defparam \a_data5[0] .power_up = "low";

dffeas \a_data3[0] (
	.clk(clk),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_data3[0]~q ),
	.prn(vcc));
defparam \a_data3[0] .is_wysiwyg = "true";
defparam \a_data3[0] .power_up = "low";

dffeas \a_data1[0] (
	.clk(clk),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_data1[0]~q ),
	.prn(vcc));
defparam \a_data1[0] .is_wysiwyg = "true";
defparam \a_data1[0] .power_up = "low";

cycloneive_lcell_comb \Mux1~0 (
	.dataa(state_register_1),
	.datab(\a_data3[0]~q ),
	.datac(state_register_0),
	.datad(\a_data1[0]~q ),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hE5E0;
defparam \Mux1~0 .sum_lutc_input = "datac";

dffeas \a_data7[0] (
	.clk(clk),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_data7[0]~q ),
	.prn(vcc));
defparam \a_data7[0] .is_wysiwyg = "true";
defparam \a_data7[0] .power_up = "low";

cycloneive_lcell_comb \Mux1~1 (
	.dataa(\a_data5[0]~q ),
	.datab(state_register_1),
	.datac(\Mux1~0_combout ),
	.datad(\a_data7[0]~q ),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
defparam \Mux1~1 .lut_mask = 16'hF838;
defparam \Mux1~1 .sum_lutc_input = "datac";

dffeas \a_channel[2] (
	.clk(clk),
	.d(in_channel[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_channel[2]~q ),
	.prn(vcc));
defparam \a_channel[2] .is_wysiwyg = "true";
defparam \a_channel[2] .power_up = "low";

dffeas \a_channel[1] (
	.clk(clk),
	.d(in_channel[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_channel[1]~q ),
	.prn(vcc));
defparam \a_channel[1] .is_wysiwyg = "true";
defparam \a_channel[1] .power_up = "low";

dffeas \a_channel[0] (
	.clk(clk),
	.d(in_channel[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_channel[0]~q ),
	.prn(vcc));
defparam \a_channel[0] .is_wysiwyg = "true";
defparam \a_channel[0] .power_up = "low";

dffeas \a_channel[8] (
	.clk(clk),
	.d(in_channel[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_channel[8]~q ),
	.prn(vcc));
defparam \a_channel[8] .is_wysiwyg = "true";
defparam \a_channel[8] .power_up = "low";

endmodule

module flashLoader_adapter_8_4 (
	reset_n,
	in_channel,
	out_valid1,
	request_1,
	full_addercout_1,
	cout,
	mem_used_9,
	request_2,
	cout1,
	state_register_0,
	always4,
	always41,
	a_valid1,
	in_ready1,
	out_endofpacket1,
	in_valid,
	out_data_0,
	out_channel_2,
	out_channel_1,
	out_channel_0,
	out_channel_8,
	in_endofpacket,
	in_data,
	clk)/* synthesis synthesis_greybox=0 */;
input 	reset_n;
input 	[11:0] in_channel;
output 	out_valid1;
input 	request_1;
input 	full_addercout_1;
input 	cout;
input 	mem_used_9;
input 	request_2;
input 	cout1;
output 	state_register_0;
output 	always4;
output 	always41;
output 	a_valid1;
output 	in_ready1;
output 	out_endofpacket1;
input 	in_valid;
output 	out_data_0;
output 	out_channel_2;
output 	out_channel_1;
output 	out_channel_0;
output 	out_channel_8;
input 	in_endofpacket;
input 	[7:0] in_data;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always4~2_combout ;
wire \state_register[0]~0_combout ;
wire \a_endofpacket~q ;
wire \Mux4~0_combout ;
wire \a_data7[0]~q ;
wire \a_data3[0]~q ;
wire \b_data[0]~0_combout ;
wire \a_channel[2]~q ;
wire \a_channel[1]~q ;
wire \a_channel[0]~q ;
wire \a_channel[8]~q ;


dffeas out_valid(
	.clk(clk),
	.d(a_valid1),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.q(out_valid1),
	.prn(vcc));
defparam out_valid.is_wysiwyg = "true";
defparam out_valid.power_up = "low";

dffeas \state_register[0] (
	.clk(clk),
	.d(\state_register[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(state_register_0),
	.prn(vcc));
defparam \state_register[0] .is_wysiwyg = "true";
defparam \state_register[0] .power_up = "low";

cycloneive_lcell_comb \always4~0 (
	.dataa(cout1),
	.datab(request_1),
	.datac(request_2),
	.datad(mem_used_9),
	.cin(gnd),
	.combout(always4),
	.cout());
defparam \always4~0 .lut_mask = 16'h002D;
defparam \always4~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always4~1 (
	.dataa(full_addercout_1),
	.datab(cout),
	.datac(mem_used_9),
	.datad(out_valid1),
	.cin(gnd),
	.combout(always41),
	.cout());
defparam \always4~1 .lut_mask = 16'h09FF;
defparam \always4~1 .sum_lutc_input = "datac";

dffeas a_valid(
	.clk(clk),
	.d(in_valid),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(a_valid1),
	.prn(vcc));
defparam a_valid.is_wysiwyg = "true";
defparam a_valid.power_up = "low";

cycloneive_lcell_comb in_ready(
	.dataa(state_register_0),
	.datab(always4),
	.datac(always41),
	.datad(a_valid1),
	.cin(gnd),
	.combout(in_ready1),
	.cout());
defparam in_ready.lut_mask = 16'hA8FF;
defparam in_ready.sum_lutc_input = "datac";

dffeas out_endofpacket(
	.clk(clk),
	.d(\Mux4~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.q(out_endofpacket1),
	.prn(vcc));
defparam out_endofpacket.is_wysiwyg = "true";
defparam out_endofpacket.power_up = "low";

dffeas \out_data[0] (
	.clk(clk),
	.d(\b_data[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.q(out_data_0),
	.prn(vcc));
defparam \out_data[0] .is_wysiwyg = "true";
defparam \out_data[0] .power_up = "low";

dffeas \out_channel[2] (
	.clk(clk),
	.d(\a_channel[2]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.q(out_channel_2),
	.prn(vcc));
defparam \out_channel[2] .is_wysiwyg = "true";
defparam \out_channel[2] .power_up = "low";

dffeas \out_channel[1] (
	.clk(clk),
	.d(\a_channel[1]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.q(out_channel_1),
	.prn(vcc));
defparam \out_channel[1] .is_wysiwyg = "true";
defparam \out_channel[1] .power_up = "low";

dffeas \out_channel[0] (
	.clk(clk),
	.d(\a_channel[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.q(out_channel_0),
	.prn(vcc));
defparam \out_channel[0] .is_wysiwyg = "true";
defparam \out_channel[0] .power_up = "low";

dffeas \out_channel[8] (
	.clk(clk),
	.d(\a_channel[8]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.q(out_channel_8),
	.prn(vcc));
defparam \out_channel[8] .is_wysiwyg = "true";
defparam \out_channel[8] .power_up = "low";

cycloneive_lcell_comb \always4~2 (
	.dataa(always4),
	.datab(always41),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\always4~2_combout ),
	.cout());
defparam \always4~2 .lut_mask = 16'hEEEE;
defparam \always4~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \state_register[0]~0 (
	.dataa(always4),
	.datab(always41),
	.datac(state_register_0),
	.datad(a_valid1),
	.cin(gnd),
	.combout(\state_register[0]~0_combout ),
	.cout());
defparam \state_register[0]~0 .lut_mask = 16'h1EF0;
defparam \state_register[0]~0 .sum_lutc_input = "datac";

dffeas a_endofpacket(
	.clk(clk),
	.d(in_endofpacket),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_endofpacket~q ),
	.prn(vcc));
defparam a_endofpacket.is_wysiwyg = "true";
defparam a_endofpacket.power_up = "low";

cycloneive_lcell_comb \Mux4~0 (
	.dataa(a_valid1),
	.datab(state_register_0),
	.datac(\a_endofpacket~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
defparam \Mux4~0 .lut_mask = 16'h8080;
defparam \Mux4~0 .sum_lutc_input = "datac";

dffeas \a_data7[0] (
	.clk(clk),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_data7[0]~q ),
	.prn(vcc));
defparam \a_data7[0] .is_wysiwyg = "true";
defparam \a_data7[0] .power_up = "low";

dffeas \a_data3[0] (
	.clk(clk),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_data3[0]~q ),
	.prn(vcc));
defparam \a_data3[0] .is_wysiwyg = "true";
defparam \a_data3[0] .power_up = "low";

cycloneive_lcell_comb \b_data[0]~0 (
	.dataa(\a_data7[0]~q ),
	.datab(\a_data3[0]~q ),
	.datac(gnd),
	.datad(state_register_0),
	.cin(gnd),
	.combout(\b_data[0]~0_combout ),
	.cout());
defparam \b_data[0]~0 .lut_mask = 16'hAACC;
defparam \b_data[0]~0 .sum_lutc_input = "datac";

dffeas \a_channel[2] (
	.clk(clk),
	.d(in_channel[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_channel[2]~q ),
	.prn(vcc));
defparam \a_channel[2] .is_wysiwyg = "true";
defparam \a_channel[2] .power_up = "low";

dffeas \a_channel[1] (
	.clk(clk),
	.d(in_channel[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_channel[1]~q ),
	.prn(vcc));
defparam \a_channel[1] .is_wysiwyg = "true";
defparam \a_channel[1] .power_up = "low";

dffeas \a_channel[0] (
	.clk(clk),
	.d(in_channel[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_channel[0]~q ),
	.prn(vcc));
defparam \a_channel[0] .is_wysiwyg = "true";
defparam \a_channel[0] .power_up = "low";

dffeas \a_channel[8] (
	.clk(clk),
	.d(in_channel[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_channel[8]~q ),
	.prn(vcc));
defparam \a_channel[8] .is_wysiwyg = "true";
defparam \a_channel[8] .power_up = "low";

endmodule

module flashLoader_clk_div (
	csr_clk_baud_rate_data_0,
	reset,
	csr_clk_baud_rate_data_1,
	csr_clk_baud_rate_data_2,
	csr_clk_baud_rate_data_3,
	csr_clk_baud_rate_data_4,
	stateST_DEASSERT_CS_DLY,
	WideOr7,
	clk_track1,
	clk_out,
	Equal0,
	Equal01,
	enable_d1,
	Add1,
	enable,
	Equal02,
	rising_edge1,
	clk)/* synthesis synthesis_greybox=0 */;
input 	csr_clk_baud_rate_data_0;
input 	reset;
input 	csr_clk_baud_rate_data_1;
input 	csr_clk_baud_rate_data_2;
input 	csr_clk_baud_rate_data_3;
input 	csr_clk_baud_rate_data_4;
input 	stateST_DEASSERT_CS_DLY;
input 	WideOr7;
output 	clk_track1;
output 	clk_out;
output 	Equal0;
output 	Equal01;
output 	enable_d1;
output 	Add1;
input 	enable;
output 	Equal02;
output 	rising_edge1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \clk_track~2_combout ;
wire \Add0~1 ;
wire \Add0~3 ;
wire \Add0~5 ;
wire \Add0~7 ;
wire \Add0~8_combout ;
wire \Add0~4_combout ;
wire \Add0~2_combout ;
wire \Add0~0_combout ;
wire \cnt_reg~3_combout ;
wire \cnt_reg[0]~q ;
wire \Add1~4_combout ;
wire \cnt_reg~2_combout ;
wire \cnt_reg[1]~q ;
wire \Add1~3_combout ;
wire \cnt_reg~1_combout ;
wire \cnt_reg[2]~q ;
wire \Add0~6_combout ;
wire \cnt_reg~4_combout ;
wire \cnt_reg[3]~q ;
wire \Add1~0_combout ;
wire \Add1~2_combout ;
wire \cnt_reg~0_combout ;
wire \cnt_reg[4]~q ;
wire \Equal0~0_combout ;
wire \clk_track_d~0_combout ;
wire \clk_track_d~q ;


dffeas clk_track(
	.clk(clk),
	.d(\clk_track~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(clk_track1),
	.prn(vcc));
defparam clk_track.is_wysiwyg = "true";
defparam clk_track.power_up = "low";

cycloneive_lcell_comb \clk_out~0 (
	.dataa(stateST_DEASSERT_CS_DLY),
	.datab(WideOr7),
	.datac(gnd),
	.datad(clk_track1),
	.cin(gnd),
	.combout(clk_out),
	.cout());
defparam \clk_out~0 .lut_mask = 16'hEEFF;
defparam \clk_out~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(csr_clk_baud_rate_data_4),
	.datab(\cnt_reg[4]~q ),
	.datac(\Add1~0_combout ),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(Equal0),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h0096;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(csr_clk_baud_rate_data_1),
	.datab(\cnt_reg[1]~q ),
	.datac(csr_clk_baud_rate_data_0),
	.datad(\cnt_reg[0]~q ),
	.cin(gnd),
	.combout(Equal01),
	.cout());
defparam \Equal0~2 .lut_mask = 16'h0690;
defparam \Equal0~2 .sum_lutc_input = "datac";

dffeas enable_d(
	.clk(clk),
	.d(enable),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(enable_d1),
	.prn(vcc));
defparam enable_d.is_wysiwyg = "true";
defparam enable_d.power_up = "low";

cycloneive_lcell_comb \Add1~1 (
	.dataa(\cnt_reg[3]~q ),
	.datab(\cnt_reg[2]~q ),
	.datac(\cnt_reg[1]~q ),
	.datad(\cnt_reg[0]~q ),
	.cin(gnd),
	.combout(Add1),
	.cout());
defparam \Add1~1 .lut_mask = 16'h6AAA;
defparam \Add1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~3 (
	.dataa(Equal0),
	.datab(Equal01),
	.datac(csr_clk_baud_rate_data_3),
	.datad(Add1),
	.cin(gnd),
	.combout(Equal02),
	.cout());
defparam \Equal0~3 .lut_mask = 16'h8008;
defparam \Equal0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb rising_edge(
	.dataa(gnd),
	.datab(gnd),
	.datac(clk_track1),
	.datad(\clk_track_d~q ),
	.cin(gnd),
	.combout(rising_edge1),
	.cout());
defparam rising_edge.lut_mask = 16'h000F;
defparam rising_edge.sum_lutc_input = "datac";

cycloneive_lcell_comb \clk_track~2 (
	.dataa(stateST_DEASSERT_CS_DLY),
	.datab(WideOr7),
	.datac(clk_track1),
	.datad(Equal02),
	.cin(gnd),
	.combout(\clk_track~2_combout ),
	.cout());
defparam \clk_track~2 .lut_mask = 16'h0110;
defparam \clk_track~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~0 (
	.dataa(csr_clk_baud_rate_data_0),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
defparam \Add0~0 .lut_mask = 16'h55AA;
defparam \Add0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~2 (
	.dataa(csr_clk_baud_rate_data_1),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
defparam \Add0~2 .lut_mask = 16'hA505;
defparam \Add0~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~4 (
	.dataa(csr_clk_baud_rate_data_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
defparam \Add0~4 .lut_mask = 16'h5AAF;
defparam \Add0~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~6 (
	.dataa(csr_clk_baud_rate_data_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
defparam \Add0~6 .lut_mask = 16'hA505;
defparam \Add0~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add0~8 (
	.dataa(csr_clk_baud_rate_data_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout());
defparam \Add0~8 .lut_mask = 16'hA5A5;
defparam \Add0~8 .sum_lutc_input = "cin";

cycloneive_lcell_comb \cnt_reg~3 (
	.dataa(\Add0~0_combout ),
	.datab(enable),
	.datac(\cnt_reg[0]~q ),
	.datad(Equal02),
	.cin(gnd),
	.combout(\cnt_reg~3_combout ),
	.cout());
defparam \cnt_reg~3 .lut_mask = 16'h222E;
defparam \cnt_reg~3 .sum_lutc_input = "datac";

dffeas \cnt_reg[0] (
	.clk(clk),
	.d(\cnt_reg~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\cnt_reg[0]~q ),
	.prn(vcc));
defparam \cnt_reg[0] .is_wysiwyg = "true";
defparam \cnt_reg[0] .power_up = "low";

cycloneive_lcell_comb \Add1~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\cnt_reg[1]~q ),
	.datad(\cnt_reg[0]~q ),
	.cin(gnd),
	.combout(\Add1~4_combout ),
	.cout());
defparam \Add1~4 .lut_mask = 16'h0FF0;
defparam \Add1~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cnt_reg~2 (
	.dataa(\Add0~2_combout ),
	.datab(enable),
	.datac(\Add1~4_combout ),
	.datad(Equal02),
	.cin(gnd),
	.combout(\cnt_reg~2_combout ),
	.cout());
defparam \cnt_reg~2 .lut_mask = 16'h22E2;
defparam \cnt_reg~2 .sum_lutc_input = "datac";

dffeas \cnt_reg[1] (
	.clk(clk),
	.d(\cnt_reg~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\cnt_reg[1]~q ),
	.prn(vcc));
defparam \cnt_reg[1] .is_wysiwyg = "true";
defparam \cnt_reg[1] .power_up = "low";

cycloneive_lcell_comb \Add1~3 (
	.dataa(gnd),
	.datab(\cnt_reg[2]~q ),
	.datac(\cnt_reg[1]~q ),
	.datad(\cnt_reg[0]~q ),
	.cin(gnd),
	.combout(\Add1~3_combout ),
	.cout());
defparam \Add1~3 .lut_mask = 16'h3CCC;
defparam \Add1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cnt_reg~1 (
	.dataa(\Add0~4_combout ),
	.datab(enable),
	.datac(\Add1~3_combout ),
	.datad(Equal02),
	.cin(gnd),
	.combout(\cnt_reg~1_combout ),
	.cout());
defparam \cnt_reg~1 .lut_mask = 16'h22E2;
defparam \cnt_reg~1 .sum_lutc_input = "datac";

dffeas \cnt_reg[2] (
	.clk(clk),
	.d(\cnt_reg~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\cnt_reg[2]~q ),
	.prn(vcc));
defparam \cnt_reg[2] .is_wysiwyg = "true";
defparam \cnt_reg[2] .power_up = "low";

cycloneive_lcell_comb \cnt_reg~4 (
	.dataa(\Add0~6_combout ),
	.datab(enable),
	.datac(Add1),
	.datad(Equal02),
	.cin(gnd),
	.combout(\cnt_reg~4_combout ),
	.cout());
defparam \cnt_reg~4 .lut_mask = 16'h22E2;
defparam \cnt_reg~4 .sum_lutc_input = "datac";

dffeas \cnt_reg[3] (
	.clk(clk),
	.d(\cnt_reg~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\cnt_reg[3]~q ),
	.prn(vcc));
defparam \cnt_reg[3] .is_wysiwyg = "true";
defparam \cnt_reg[3] .power_up = "low";

cycloneive_lcell_comb \Add1~0 (
	.dataa(\cnt_reg[2]~q ),
	.datab(\cnt_reg[1]~q ),
	.datac(\cnt_reg[0]~q ),
	.datad(\cnt_reg[3]~q ),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout());
defparam \Add1~0 .lut_mask = 16'h8000;
defparam \Add1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\cnt_reg[4]~q ),
	.datad(\Add1~0_combout ),
	.cin(gnd),
	.combout(\Add1~2_combout ),
	.cout());
defparam \Add1~2 .lut_mask = 16'h0FF0;
defparam \Add1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cnt_reg~0 (
	.dataa(\Add0~8_combout ),
	.datab(enable),
	.datac(\Add1~2_combout ),
	.datad(Equal02),
	.cin(gnd),
	.combout(\cnt_reg~0_combout ),
	.cout());
defparam \cnt_reg~0 .lut_mask = 16'h22E2;
defparam \cnt_reg~0 .sum_lutc_input = "datac";

dffeas \cnt_reg[4] (
	.clk(clk),
	.d(\cnt_reg~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\cnt_reg[4]~q ),
	.prn(vcc));
defparam \cnt_reg[4] .is_wysiwyg = "true";
defparam \cnt_reg[4] .power_up = "low";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\cnt_reg[1]~q ),
	.datab(\cnt_reg[0]~q ),
	.datac(csr_clk_baud_rate_data_2),
	.datad(\cnt_reg[2]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h8778;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \clk_track_d~0 (
	.dataa(clk_track1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\clk_track_d~0_combout ),
	.cout());
defparam \clk_track_d~0 .lut_mask = 16'h5555;
defparam \clk_track_d~0 .sum_lutc_input = "datac";

dffeas clk_track_d(
	.clk(clk),
	.d(\clk_track_d~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\clk_track_d~q ),
	.prn(vcc));
defparam clk_track_d.is_wysiwyg = "true";
defparam clk_track_d.power_up = "low";

endmodule

module flashLoader_demultiplexer_12_channels (
	data_num_lines_1,
	data_num_lines_2,
	addr_num_lines_2,
	addr_num_lines_1,
	in_cmd_channel_reg_1,
	in_cmd_channel_reg_0,
	op_num_lines_1,
	in_ready,
	data_num_lines_0,
	op_num_lines_0,
	state_register_1,
	state_register_0,
	a_valid,
	always4,
	WideOr0,
	state_register_01,
	always41,
	always42,
	a_valid1,
	in_ready1,
	op_num_lines_2,
	WideOr01,
	Selector8,
	demux_channel_2,
	Equal0,
	demux_channel_21,
	sink_ready,
	in_ready2,
	demux_channel_1,
	demux_channel_11,
	addr_num_lines_0,
	demux_channel_0,
	demux_channel_01,
	WideOr02,
	WideOr03,
	WideOr04,
	WideOr05,
	demux_channel_22,
	src0_valid1,
	src1_valid1,
	src2_valid1,
	WideOr06)/* synthesis synthesis_greybox=0 */;
input 	data_num_lines_1;
input 	data_num_lines_2;
input 	addr_num_lines_2;
input 	addr_num_lines_1;
input 	in_cmd_channel_reg_1;
input 	in_cmd_channel_reg_0;
input 	op_num_lines_1;
input 	in_ready;
input 	data_num_lines_0;
input 	op_num_lines_0;
input 	state_register_1;
input 	state_register_0;
input 	a_valid;
input 	always4;
output 	WideOr0;
input 	state_register_01;
input 	always41;
input 	always42;
input 	a_valid1;
input 	in_ready1;
input 	op_num_lines_2;
output 	WideOr01;
input 	Selector8;
input 	demux_channel_2;
input 	Equal0;
input 	demux_channel_21;
output 	sink_ready;
input 	in_ready2;
input 	demux_channel_1;
input 	demux_channel_11;
input 	addr_num_lines_0;
input 	demux_channel_0;
input 	demux_channel_01;
output 	WideOr02;
output 	WideOr03;
output 	WideOr04;
output 	WideOr05;
input 	demux_channel_22;
output 	src0_valid1;
output 	src1_valid1;
output 	src2_valid1;
output 	WideOr06;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \WideOr0~0_combout ;
wire \WideOr0~1_combout ;
wire \WideOr0~2_combout ;
wire \WideOr0~6_combout ;
wire \WideOr0~9_combout ;
wire \WideOr0~10_combout ;
wire \WideOr0~12_combout ;


cycloneive_lcell_comb \WideOr0~3 (
	.dataa(\WideOr0~0_combout ),
	.datab(in_ready),
	.datac(\WideOr0~1_combout ),
	.datad(\WideOr0~2_combout ),
	.cin(gnd),
	.combout(WideOr0),
	.cout());
defparam \WideOr0~3 .lut_mask = 16'hC0EA;
defparam \WideOr0~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~4 (
	.dataa(data_num_lines_2),
	.datab(op_num_lines_2),
	.datac(in_cmd_channel_reg_1),
	.datad(in_cmd_channel_reg_0),
	.cin(gnd),
	.combout(WideOr01),
	.cout());
defparam \WideOr0~4 .lut_mask = 16'hAACA;
defparam \WideOr0~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sink_ready~0 (
	.dataa(in_ready1),
	.datab(demux_channel_21),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(sink_ready),
	.cout());
defparam \sink_ready~0 .lut_mask = 16'h8888;
defparam \sink_ready~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~5 (
	.dataa(in_ready),
	.datab(in_ready2),
	.datac(demux_channel_11),
	.datad(demux_channel_01),
	.cin(gnd),
	.combout(WideOr02),
	.cout());
defparam \WideOr0~5 .lut_mask = 16'hEAC0;
defparam \WideOr0~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~7 (
	.dataa(WideOr01),
	.datab(state_register_01),
	.datac(always41),
	.datad(\WideOr0~6_combout ),
	.cin(gnd),
	.combout(WideOr03),
	.cout());
defparam \WideOr0~7 .lut_mask = 16'hAA80;
defparam \WideOr0~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~8 (
	.dataa(in_ready),
	.datab(in_ready2),
	.datac(op_num_lines_1),
	.datad(op_num_lines_0),
	.cin(gnd),
	.combout(WideOr04),
	.cout());
defparam \WideOr0~8 .lut_mask = 16'hEAC0;
defparam \WideOr0~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~11 (
	.dataa(Equal0),
	.datab(WideOr04),
	.datac(\WideOr0~9_combout ),
	.datad(\WideOr0~10_combout ),
	.cin(gnd),
	.combout(WideOr05),
	.cout());
defparam \WideOr0~11 .lut_mask = 16'hFDF8;
defparam \WideOr0~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb src0_valid(
	.dataa(Selector8),
	.datab(op_num_lines_0),
	.datac(demux_channel_0),
	.datad(demux_channel_22),
	.cin(gnd),
	.combout(src0_valid1),
	.cout());
defparam src0_valid.lut_mask = 16'h88A0;
defparam src0_valid.sum_lutc_input = "datac";

cycloneive_lcell_comb src1_valid(
	.dataa(Selector8),
	.datab(op_num_lines_1),
	.datac(demux_channel_1),
	.datad(demux_channel_22),
	.cin(gnd),
	.combout(src1_valid1),
	.cout());
defparam src1_valid.lut_mask = 16'h88A0;
defparam src1_valid.sum_lutc_input = "datac";

cycloneive_lcell_comb src2_valid(
	.dataa(Selector8),
	.datab(op_num_lines_2),
	.datac(demux_channel_2),
	.datad(demux_channel_22),
	.cin(gnd),
	.combout(src2_valid1),
	.cout());
defparam src2_valid.lut_mask = 16'h88A0;
defparam src2_valid.sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~13 (
	.dataa(in_ready2),
	.datab(op_num_lines_1),
	.datac(\WideOr0~12_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(WideOr06),
	.cout());
defparam \WideOr0~13 .lut_mask = 16'hF8F8;
defparam \WideOr0~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~0 (
	.dataa(data_num_lines_1),
	.datab(op_num_lines_1),
	.datac(in_cmd_channel_reg_1),
	.datad(in_cmd_channel_reg_0),
	.cin(gnd),
	.combout(\WideOr0~0_combout ),
	.cout());
defparam \WideOr0~0 .lut_mask = 16'hAACA;
defparam \WideOr0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~1 (
	.dataa(in_cmd_channel_reg_1),
	.datab(in_cmd_channel_reg_0),
	.datac(data_num_lines_0),
	.datad(op_num_lines_0),
	.cin(gnd),
	.combout(\WideOr0~1_combout ),
	.cout());
defparam \WideOr0~1 .lut_mask = 16'hF2D0;
defparam \WideOr0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~2 (
	.dataa(state_register_1),
	.datab(state_register_0),
	.datac(a_valid),
	.datad(always4),
	.cin(gnd),
	.combout(\WideOr0~2_combout ),
	.cout());
defparam \WideOr0~2 .lut_mask = 16'h70F0;
defparam \WideOr0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~6 (
	.dataa(state_register_01),
	.datab(always42),
	.datac(a_valid1),
	.datad(gnd),
	.cin(gnd),
	.combout(\WideOr0~6_combout ),
	.cout());
defparam \WideOr0~6 .lut_mask = 16'h8F8F;
defparam \WideOr0~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~9 (
	.dataa(Equal0),
	.datab(in_ready1),
	.datac(op_num_lines_2),
	.datad(addr_num_lines_2),
	.cin(gnd),
	.combout(\WideOr0~9_combout ),
	.cout());
defparam \WideOr0~9 .lut_mask = 16'hC480;
defparam \WideOr0~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~10 (
	.dataa(in_ready),
	.datab(addr_num_lines_0),
	.datac(in_ready2),
	.datad(addr_num_lines_1),
	.cin(gnd),
	.combout(\WideOr0~10_combout ),
	.cout());
defparam \WideOr0~10 .lut_mask = 16'hF888;
defparam \WideOr0~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr0~12 (
	.dataa(in_ready1),
	.datab(op_num_lines_2),
	.datac(in_ready),
	.datad(op_num_lines_0),
	.cin(gnd),
	.combout(\WideOr0~12_combout ),
	.cout());
defparam \WideOr0~12 .lut_mask = 16'hF888;
defparam \WideOr0~12 .sum_lutc_input = "datac";

endmodule

module flashLoader_inf_sc_fifo_ser_data (
	altera_reset_synchronizer_int_chain_out,
	out_payload_12,
	out_payload_2,
	out_payload_1,
	out_payload_0,
	mem_used_9,
	out_valid,
	stateST_SEND,
	fifo_pop_out,
	out_payload_16,
	out_payload_8,
	WideOr1,
	write,
	src_payload_0,
	src_data_0,
	src_channel_2,
	src_channel_1,
	src_channel_0,
	src_channel_8,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	altera_reset_synchronizer_int_chain_out;
output 	out_payload_12;
output 	out_payload_2;
output 	out_payload_1;
output 	out_payload_0;
output 	mem_used_9;
output 	out_valid;
input 	stateST_SEND;
input 	fifo_pop_out;
output 	out_payload_16;
output 	out_payload_8;
input 	WideOr1;
output 	write;
input 	src_payload_0;
input 	src_data_0;
input 	src_channel_2;
input 	src_channel_1;
input 	src_channel_0;
input 	src_channel_8;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



flashLoader_altera_avalon_sc_fifo inf_sc_fifo_ser_data(
	.reset(altera_reset_synchronizer_int_chain_out),
	.out_payload_12(out_payload_12),
	.out_payload_2(out_payload_2),
	.out_payload_1(out_payload_1),
	.out_payload_0(out_payload_0),
	.mem_used_9(mem_used_9),
	.out_valid1(out_valid),
	.stateST_SEND(stateST_SEND),
	.fifo_pop_out(fifo_pop_out),
	.out_payload_16(out_payload_16),
	.out_payload_8(out_payload_8),
	.WideOr1(WideOr1),
	.write(write),
	.src_payload_0(src_payload_0),
	.src_data_0(src_data_0),
	.src_channel_2(src_channel_2),
	.src_channel_1(src_channel_1),
	.src_channel_0(src_channel_0),
	.src_channel_8(src_channel_8),
	.clk(clk_clk));

endmodule

module flashLoader_altera_avalon_sc_fifo (
	reset,
	out_payload_12,
	out_payload_2,
	out_payload_1,
	out_payload_0,
	mem_used_9,
	out_valid1,
	stateST_SEND,
	fifo_pop_out,
	out_payload_16,
	out_payload_8,
	WideOr1,
	write,
	src_payload_0,
	src_data_0,
	src_channel_2,
	src_channel_1,
	src_channel_0,
	src_channel_8,
	clk)/* synthesis synthesis_greybox=0 */;
input 	reset;
output 	out_payload_12;
output 	out_payload_2;
output 	out_payload_1;
output 	out_payload_0;
output 	mem_used_9;
output 	out_valid1;
input 	stateST_SEND;
input 	fifo_pop_out;
output 	out_payload_16;
output 	out_payload_8;
input 	WideOr1;
output 	write;
input 	src_payload_0;
input 	src_data_0;
input 	src_channel_2;
input 	src_channel_1;
input 	src_channel_0;
input 	src_channel_8;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem[9][12]~q ;
wire \mem~48_combout ;
wire \internal_out_ready~combout ;
wire \read~0_combout ;
wire \mem_used~1_combout ;
wire \mem_used[8]~2_combout ;
wire \mem_used[8]~q ;
wire \mem_used~5_combout ;
wire \mem_used[7]~q ;
wire \mem_used~7_combout ;
wire \mem_used[6]~q ;
wire \mem_used~9_combout ;
wire \mem_used[5]~q ;
wire \mem_used~10_combout ;
wire \mem_used[4]~q ;
wire \mem_used~8_combout ;
wire \mem_used[3]~q ;
wire \mem_used~6_combout ;
wire \mem_used[2]~q ;
wire \mem_used~3_combout ;
wire \mem_used[1]~q ;
wire \mem_used[0]~4_combout ;
wire \mem_used[0]~q ;
wire \internal_out_valid~0_combout ;
wire \internal_out_valid~q ;
wire \always8~0_combout ;
wire \mem[8][12]~q ;
wire \mem~42_combout ;
wire \always7~0_combout ;
wire \mem[7][12]~q ;
wire \mem~36_combout ;
wire \always6~0_combout ;
wire \mem[6][12]~q ;
wire \mem~30_combout ;
wire \always5~0_combout ;
wire \mem[5][12]~q ;
wire \mem~24_combout ;
wire \always4~0_combout ;
wire \mem[4][12]~q ;
wire \mem~18_combout ;
wire \always3~0_combout ;
wire \mem[3][12]~q ;
wire \mem~12_combout ;
wire \always2~0_combout ;
wire \mem[2][12]~q ;
wire \mem~6_combout ;
wire \always1~0_combout ;
wire \mem[1][12]~q ;
wire \mem~0_combout ;
wire \mem[0][12]~q ;
wire \mem[9][2]~q ;
wire \mem~49_combout ;
wire \mem[8][2]~q ;
wire \mem~43_combout ;
wire \mem[7][2]~q ;
wire \mem~37_combout ;
wire \mem[6][2]~q ;
wire \mem~31_combout ;
wire \mem[5][2]~q ;
wire \mem~25_combout ;
wire \mem[4][2]~q ;
wire \mem~19_combout ;
wire \mem[3][2]~q ;
wire \mem~13_combout ;
wire \mem[2][2]~q ;
wire \mem~7_combout ;
wire \mem[1][2]~q ;
wire \mem~1_combout ;
wire \mem[0][2]~q ;
wire \mem[9][1]~q ;
wire \mem~50_combout ;
wire \mem[8][1]~q ;
wire \mem~44_combout ;
wire \mem[7][1]~q ;
wire \mem~38_combout ;
wire \mem[6][1]~q ;
wire \mem~32_combout ;
wire \mem[5][1]~q ;
wire \mem~26_combout ;
wire \mem[4][1]~q ;
wire \mem~20_combout ;
wire \mem[3][1]~q ;
wire \mem~14_combout ;
wire \mem[2][1]~q ;
wire \mem~8_combout ;
wire \mem[1][1]~q ;
wire \mem~2_combout ;
wire \mem[0][1]~q ;
wire \mem[9][0]~q ;
wire \mem~51_combout ;
wire \mem[8][0]~q ;
wire \mem~45_combout ;
wire \mem[7][0]~q ;
wire \mem~39_combout ;
wire \mem[6][0]~q ;
wire \mem~33_combout ;
wire \mem[5][0]~q ;
wire \mem~27_combout ;
wire \mem[4][0]~q ;
wire \mem~21_combout ;
wire \mem[3][0]~q ;
wire \mem~15_combout ;
wire \mem[2][0]~q ;
wire \mem~9_combout ;
wire \mem[1][0]~q ;
wire \mem~3_combout ;
wire \mem[0][0]~q ;
wire \mem_used[9]~0_combout ;
wire \mem[9][16]~q ;
wire \mem~52_combout ;
wire \mem[8][16]~q ;
wire \mem~46_combout ;
wire \mem[7][16]~q ;
wire \mem~40_combout ;
wire \mem[6][16]~q ;
wire \mem~34_combout ;
wire \mem[5][16]~q ;
wire \mem~28_combout ;
wire \mem[4][16]~q ;
wire \mem~22_combout ;
wire \mem[3][16]~q ;
wire \mem~16_combout ;
wire \mem[2][16]~q ;
wire \mem~10_combout ;
wire \mem[1][16]~q ;
wire \mem~4_combout ;
wire \mem[0][16]~q ;
wire \mem[9][8]~q ;
wire \mem~53_combout ;
wire \mem[8][8]~q ;
wire \mem~47_combout ;
wire \mem[7][8]~q ;
wire \mem~41_combout ;
wire \mem[6][8]~q ;
wire \mem~35_combout ;
wire \mem[5][8]~q ;
wire \mem~29_combout ;
wire \mem[4][8]~q ;
wire \mem~23_combout ;
wire \mem[3][8]~q ;
wire \mem~17_combout ;
wire \mem[2][8]~q ;
wire \mem~11_combout ;
wire \mem[1][8]~q ;
wire \mem~5_combout ;
wire \mem[0][8]~q ;


dffeas \out_payload[12] (
	.clk(clk),
	.d(\mem[0][12]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_12),
	.prn(vcc));
defparam \out_payload[12] .is_wysiwyg = "true";
defparam \out_payload[12] .power_up = "low";

dffeas \out_payload[2] (
	.clk(clk),
	.d(\mem[0][2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_2),
	.prn(vcc));
defparam \out_payload[2] .is_wysiwyg = "true";
defparam \out_payload[2] .power_up = "low";

dffeas \out_payload[1] (
	.clk(clk),
	.d(\mem[0][1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_1),
	.prn(vcc));
defparam \out_payload[1] .is_wysiwyg = "true";
defparam \out_payload[1] .power_up = "low";

dffeas \out_payload[0] (
	.clk(clk),
	.d(\mem[0][0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_0),
	.prn(vcc));
defparam \out_payload[0] .is_wysiwyg = "true";
defparam \out_payload[0] .power_up = "low";

dffeas \mem_used[9] (
	.clk(clk),
	.d(\mem_used[9]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_9),
	.prn(vcc));
defparam \mem_used[9] .is_wysiwyg = "true";
defparam \mem_used[9] .power_up = "low";

dffeas out_valid(
	.clk(clk),
	.d(\internal_out_valid~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_valid1),
	.prn(vcc));
defparam out_valid.is_wysiwyg = "true";
defparam out_valid.power_up = "low";

dffeas \out_payload[16] (
	.clk(clk),
	.d(\mem[0][16]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_16),
	.prn(vcc));
defparam \out_payload[16] .is_wysiwyg = "true";
defparam \out_payload[16] .power_up = "low";

dffeas \out_payload[8] (
	.clk(clk),
	.d(\mem[0][8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_8),
	.prn(vcc));
defparam \out_payload[8] .is_wysiwyg = "true";
defparam \out_payload[8] .power_up = "low";

cycloneive_lcell_comb \write~0 (
	.dataa(WideOr1),
	.datab(gnd),
	.datac(gnd),
	.datad(mem_used_9),
	.cin(gnd),
	.combout(write),
	.cout());
defparam \write~0 .lut_mask = 16'h00AA;
defparam \write~0 .sum_lutc_input = "datac";

dffeas \mem[9][12] (
	.clk(clk),
	.d(\mem~48_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[9][12]~q ),
	.prn(vcc));
defparam \mem[9][12] .is_wysiwyg = "true";
defparam \mem[9][12] .power_up = "low";

cycloneive_lcell_comb \mem~48 (
	.dataa(\mem[9][12]~q ),
	.datab(src_data_0),
	.datac(gnd),
	.datad(mem_used_9),
	.cin(gnd),
	.combout(\mem~48_combout ),
	.cout());
defparam \mem~48 .lut_mask = 16'hAACC;
defparam \mem~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb internal_out_ready(
	.dataa(stateST_SEND),
	.datab(fifo_pop_out),
	.datac(gnd),
	.datad(out_valid1),
	.cin(gnd),
	.combout(\internal_out_ready~combout ),
	.cout());
defparam internal_out_ready.lut_mask = 16'h88FF;
defparam internal_out_ready.sum_lutc_input = "datac";

cycloneive_lcell_comb \read~0 (
	.dataa(out_valid1),
	.datab(stateST_SEND),
	.datac(fifo_pop_out),
	.datad(\internal_out_valid~q ),
	.cin(gnd),
	.combout(\read~0_combout ),
	.cout());
defparam \read~0 .lut_mask = 16'h2AFF;
defparam \read~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used~1 (
	.dataa(mem_used_9),
	.datab(WideOr1),
	.datac(\mem_used[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used~1_combout ),
	.cout());
defparam \mem_used~1 .lut_mask = 16'hEAEA;
defparam \mem_used~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_used[8]~2 (
	.dataa(WideOr1),
	.datab(mem_used_9),
	.datac(\internal_out_ready~combout ),
	.datad(\internal_out_valid~q ),
	.cin(gnd),
	.combout(\mem_used[8]~2_combout ),
	.cout());
defparam \mem_used[8]~2 .lut_mask = 16'hD222;
defparam \mem_used[8]~2 .sum_lutc_input = "datac";

dffeas \mem_used[8] (
	.clk(clk),
	.d(\mem_used~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[8]~2_combout ),
	.q(\mem_used[8]~q ),
	.prn(vcc));
defparam \mem_used[8] .is_wysiwyg = "true";
defparam \mem_used[8] .power_up = "low";

cycloneive_lcell_comb \mem_used~5 (
	.dataa(\mem_used[8]~q ),
	.datab(\mem_used[6]~q ),
	.datac(WideOr1),
	.datad(mem_used_9),
	.cin(gnd),
	.combout(\mem_used~5_combout ),
	.cout());
defparam \mem_used~5 .lut_mask = 16'hAACA;
defparam \mem_used~5 .sum_lutc_input = "datac";

dffeas \mem_used[7] (
	.clk(clk),
	.d(\mem_used~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[8]~2_combout ),
	.q(\mem_used[7]~q ),
	.prn(vcc));
defparam \mem_used[7] .is_wysiwyg = "true";
defparam \mem_used[7] .power_up = "low";

cycloneive_lcell_comb \mem_used~7 (
	.dataa(\mem_used[7]~q ),
	.datab(\mem_used[5]~q ),
	.datac(WideOr1),
	.datad(mem_used_9),
	.cin(gnd),
	.combout(\mem_used~7_combout ),
	.cout());
defparam \mem_used~7 .lut_mask = 16'hAACA;
defparam \mem_used~7 .sum_lutc_input = "datac";

dffeas \mem_used[6] (
	.clk(clk),
	.d(\mem_used~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[8]~2_combout ),
	.q(\mem_used[6]~q ),
	.prn(vcc));
defparam \mem_used[6] .is_wysiwyg = "true";
defparam \mem_used[6] .power_up = "low";

cycloneive_lcell_comb \mem_used~9 (
	.dataa(\mem_used[6]~q ),
	.datab(\mem_used[4]~q ),
	.datac(WideOr1),
	.datad(mem_used_9),
	.cin(gnd),
	.combout(\mem_used~9_combout ),
	.cout());
defparam \mem_used~9 .lut_mask = 16'hAACA;
defparam \mem_used~9 .sum_lutc_input = "datac";

dffeas \mem_used[5] (
	.clk(clk),
	.d(\mem_used~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[8]~2_combout ),
	.q(\mem_used[5]~q ),
	.prn(vcc));
defparam \mem_used[5] .is_wysiwyg = "true";
defparam \mem_used[5] .power_up = "low";

cycloneive_lcell_comb \mem_used~10 (
	.dataa(\mem_used[5]~q ),
	.datab(\mem_used[3]~q ),
	.datac(WideOr1),
	.datad(mem_used_9),
	.cin(gnd),
	.combout(\mem_used~10_combout ),
	.cout());
defparam \mem_used~10 .lut_mask = 16'hAACA;
defparam \mem_used~10 .sum_lutc_input = "datac";

dffeas \mem_used[4] (
	.clk(clk),
	.d(\mem_used~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[8]~2_combout ),
	.q(\mem_used[4]~q ),
	.prn(vcc));
defparam \mem_used[4] .is_wysiwyg = "true";
defparam \mem_used[4] .power_up = "low";

cycloneive_lcell_comb \mem_used~8 (
	.dataa(\mem_used[4]~q ),
	.datab(\mem_used[2]~q ),
	.datac(WideOr1),
	.datad(mem_used_9),
	.cin(gnd),
	.combout(\mem_used~8_combout ),
	.cout());
defparam \mem_used~8 .lut_mask = 16'hAACA;
defparam \mem_used~8 .sum_lutc_input = "datac";

dffeas \mem_used[3] (
	.clk(clk),
	.d(\mem_used~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[8]~2_combout ),
	.q(\mem_used[3]~q ),
	.prn(vcc));
defparam \mem_used[3] .is_wysiwyg = "true";
defparam \mem_used[3] .power_up = "low";

cycloneive_lcell_comb \mem_used~6 (
	.dataa(\mem_used[3]~q ),
	.datab(\mem_used[1]~q ),
	.datac(WideOr1),
	.datad(mem_used_9),
	.cin(gnd),
	.combout(\mem_used~6_combout ),
	.cout());
defparam \mem_used~6 .lut_mask = 16'hAACA;
defparam \mem_used~6 .sum_lutc_input = "datac";

dffeas \mem_used[2] (
	.clk(clk),
	.d(\mem_used~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[8]~2_combout ),
	.q(\mem_used[2]~q ),
	.prn(vcc));
defparam \mem_used[2] .is_wysiwyg = "true";
defparam \mem_used[2] .power_up = "low";

cycloneive_lcell_comb \mem_used~3 (
	.dataa(\mem_used[2]~q ),
	.datab(\mem_used[0]~q ),
	.datac(WideOr1),
	.datad(mem_used_9),
	.cin(gnd),
	.combout(\mem_used~3_combout ),
	.cout());
defparam \mem_used~3 .lut_mask = 16'hAACA;
defparam \mem_used~3 .sum_lutc_input = "datac";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[8]~2_combout ),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cycloneive_lcell_comb \mem_used[0]~4 (
	.dataa(\mem_used[0]~q ),
	.datab(write),
	.datac(\read~0_combout ),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem_used[0]~4_combout ),
	.cout());
defparam \mem_used[0]~4 .lut_mask = 16'hEBE8;
defparam \mem_used[0]~4 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cycloneive_lcell_comb \internal_out_valid~0 (
	.dataa(\mem_used[0]~q ),
	.datab(gnd),
	.datac(\internal_out_ready~combout ),
	.datad(\internal_out_valid~q ),
	.cin(gnd),
	.combout(\internal_out_valid~0_combout ),
	.cout());
defparam \internal_out_valid~0 .lut_mask = 16'h0AAA;
defparam \internal_out_valid~0 .sum_lutc_input = "datac";

dffeas internal_out_valid(
	.clk(clk),
	.d(\internal_out_valid~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_valid~q ),
	.prn(vcc));
defparam internal_out_valid.is_wysiwyg = "true";
defparam internal_out_valid.power_up = "low";

cycloneive_lcell_comb \always8~0 (
	.dataa(\internal_out_ready~combout ),
	.datab(\internal_out_valid~q ),
	.datac(gnd),
	.datad(\mem_used[8]~q ),
	.cin(gnd),
	.combout(\always8~0_combout ),
	.cout());
defparam \always8~0 .lut_mask = 16'h88FF;
defparam \always8~0 .sum_lutc_input = "datac";

dffeas \mem[8][12] (
	.clk(clk),
	.d(\mem~48_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always8~0_combout ),
	.q(\mem[8][12]~q ),
	.prn(vcc));
defparam \mem[8][12] .is_wysiwyg = "true";
defparam \mem[8][12] .power_up = "low";

cycloneive_lcell_comb \mem~42 (
	.dataa(\mem[8][12]~q ),
	.datab(src_data_0),
	.datac(gnd),
	.datad(\mem_used[8]~q ),
	.cin(gnd),
	.combout(\mem~42_combout ),
	.cout());
defparam \mem~42 .lut_mask = 16'hAACC;
defparam \mem~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always7~0 (
	.dataa(\internal_out_ready~combout ),
	.datab(\internal_out_valid~q ),
	.datac(gnd),
	.datad(\mem_used[7]~q ),
	.cin(gnd),
	.combout(\always7~0_combout ),
	.cout());
defparam \always7~0 .lut_mask = 16'h88FF;
defparam \always7~0 .sum_lutc_input = "datac";

dffeas \mem[7][12] (
	.clk(clk),
	.d(\mem~42_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\mem[7][12]~q ),
	.prn(vcc));
defparam \mem[7][12] .is_wysiwyg = "true";
defparam \mem[7][12] .power_up = "low";

cycloneive_lcell_comb \mem~36 (
	.dataa(\mem[7][12]~q ),
	.datab(src_data_0),
	.datac(gnd),
	.datad(\mem_used[7]~q ),
	.cin(gnd),
	.combout(\mem~36_combout ),
	.cout());
defparam \mem~36 .lut_mask = 16'hAACC;
defparam \mem~36 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always6~0 (
	.dataa(\internal_out_ready~combout ),
	.datab(\internal_out_valid~q ),
	.datac(gnd),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\always6~0_combout ),
	.cout());
defparam \always6~0 .lut_mask = 16'h88FF;
defparam \always6~0 .sum_lutc_input = "datac";

dffeas \mem[6][12] (
	.clk(clk),
	.d(\mem~36_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][12]~q ),
	.prn(vcc));
defparam \mem[6][12] .is_wysiwyg = "true";
defparam \mem[6][12] .power_up = "low";

cycloneive_lcell_comb \mem~30 (
	.dataa(\mem[6][12]~q ),
	.datab(src_data_0),
	.datac(gnd),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\mem~30_combout ),
	.cout());
defparam \mem~30 .lut_mask = 16'hAACC;
defparam \mem~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always5~0 (
	.dataa(\internal_out_ready~combout ),
	.datab(\internal_out_valid~q ),
	.datac(gnd),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\always5~0_combout ),
	.cout());
defparam \always5~0 .lut_mask = 16'h88FF;
defparam \always5~0 .sum_lutc_input = "datac";

dffeas \mem[5][12] (
	.clk(clk),
	.d(\mem~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\mem[5][12]~q ),
	.prn(vcc));
defparam \mem[5][12] .is_wysiwyg = "true";
defparam \mem[5][12] .power_up = "low";

cycloneive_lcell_comb \mem~24 (
	.dataa(\mem[5][12]~q ),
	.datab(src_data_0),
	.datac(gnd),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\mem~24_combout ),
	.cout());
defparam \mem~24 .lut_mask = 16'hAACC;
defparam \mem~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always4~0 (
	.dataa(\internal_out_ready~combout ),
	.datab(\internal_out_valid~q ),
	.datac(gnd),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\always4~0_combout ),
	.cout());
defparam \always4~0 .lut_mask = 16'h88FF;
defparam \always4~0 .sum_lutc_input = "datac";

dffeas \mem[4][12] (
	.clk(clk),
	.d(\mem~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(\mem[4][12]~q ),
	.prn(vcc));
defparam \mem[4][12] .is_wysiwyg = "true";
defparam \mem[4][12] .power_up = "low";

cycloneive_lcell_comb \mem~18 (
	.dataa(\mem[4][12]~q ),
	.datab(src_data_0),
	.datac(gnd),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\mem~18_combout ),
	.cout());
defparam \mem~18 .lut_mask = 16'hAACC;
defparam \mem~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always3~0 (
	.dataa(\internal_out_ready~combout ),
	.datab(\internal_out_valid~q ),
	.datac(gnd),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\always3~0_combout ),
	.cout());
defparam \always3~0 .lut_mask = 16'h88FF;
defparam \always3~0 .sum_lutc_input = "datac";

dffeas \mem[3][12] (
	.clk(clk),
	.d(\mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\mem[3][12]~q ),
	.prn(vcc));
defparam \mem[3][12] .is_wysiwyg = "true";
defparam \mem[3][12] .power_up = "low";

cycloneive_lcell_comb \mem~12 (
	.dataa(\mem[3][12]~q ),
	.datab(src_data_0),
	.datac(gnd),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\mem~12_combout ),
	.cout());
defparam \mem~12 .lut_mask = 16'hAACC;
defparam \mem~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always2~0 (
	.dataa(\internal_out_ready~combout ),
	.datab(\internal_out_valid~q ),
	.datac(gnd),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\always2~0_combout ),
	.cout());
defparam \always2~0 .lut_mask = 16'h88FF;
defparam \always2~0 .sum_lutc_input = "datac";

dffeas \mem[2][12] (
	.clk(clk),
	.d(\mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(\mem[2][12]~q ),
	.prn(vcc));
defparam \mem[2][12] .is_wysiwyg = "true";
defparam \mem[2][12] .power_up = "low";

cycloneive_lcell_comb \mem~6 (
	.dataa(\mem[2][12]~q ),
	.datab(src_data_0),
	.datac(gnd),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\mem~6_combout ),
	.cout());
defparam \mem~6 .lut_mask = 16'hAACC;
defparam \mem~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always1~0 (
	.dataa(\internal_out_ready~combout ),
	.datab(\internal_out_valid~q ),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\always1~0_combout ),
	.cout());
defparam \always1~0 .lut_mask = 16'h88FF;
defparam \always1~0 .sum_lutc_input = "datac";

dffeas \mem[1][12] (
	.clk(clk),
	.d(\mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\mem[1][12]~q ),
	.prn(vcc));
defparam \mem[1][12] .is_wysiwyg = "true";
defparam \mem[1][12] .power_up = "low";

cycloneive_lcell_comb \mem~0 (
	.dataa(\mem[1][12]~q ),
	.datab(src_data_0),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hAACC;
defparam \mem~0 .sum_lutc_input = "datac";

dffeas \mem[0][12] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\internal_out_valid~0_combout ),
	.q(\mem[0][12]~q ),
	.prn(vcc));
defparam \mem[0][12] .is_wysiwyg = "true";
defparam \mem[0][12] .power_up = "low";

dffeas \mem[9][2] (
	.clk(clk),
	.d(\mem~49_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[9][2]~q ),
	.prn(vcc));
defparam \mem[9][2] .is_wysiwyg = "true";
defparam \mem[9][2] .power_up = "low";

cycloneive_lcell_comb \mem~49 (
	.dataa(\mem[9][2]~q ),
	.datab(src_channel_2),
	.datac(gnd),
	.datad(mem_used_9),
	.cin(gnd),
	.combout(\mem~49_combout ),
	.cout());
defparam \mem~49 .lut_mask = 16'hAACC;
defparam \mem~49 .sum_lutc_input = "datac";

dffeas \mem[8][2] (
	.clk(clk),
	.d(\mem~49_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always8~0_combout ),
	.q(\mem[8][2]~q ),
	.prn(vcc));
defparam \mem[8][2] .is_wysiwyg = "true";
defparam \mem[8][2] .power_up = "low";

cycloneive_lcell_comb \mem~43 (
	.dataa(\mem[8][2]~q ),
	.datab(src_channel_2),
	.datac(gnd),
	.datad(\mem_used[8]~q ),
	.cin(gnd),
	.combout(\mem~43_combout ),
	.cout());
defparam \mem~43 .lut_mask = 16'hAACC;
defparam \mem~43 .sum_lutc_input = "datac";

dffeas \mem[7][2] (
	.clk(clk),
	.d(\mem~43_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\mem[7][2]~q ),
	.prn(vcc));
defparam \mem[7][2] .is_wysiwyg = "true";
defparam \mem[7][2] .power_up = "low";

cycloneive_lcell_comb \mem~37 (
	.dataa(\mem[7][2]~q ),
	.datab(src_channel_2),
	.datac(gnd),
	.datad(\mem_used[7]~q ),
	.cin(gnd),
	.combout(\mem~37_combout ),
	.cout());
defparam \mem~37 .lut_mask = 16'hAACC;
defparam \mem~37 .sum_lutc_input = "datac";

dffeas \mem[6][2] (
	.clk(clk),
	.d(\mem~37_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][2]~q ),
	.prn(vcc));
defparam \mem[6][2] .is_wysiwyg = "true";
defparam \mem[6][2] .power_up = "low";

cycloneive_lcell_comb \mem~31 (
	.dataa(\mem[6][2]~q ),
	.datab(src_channel_2),
	.datac(gnd),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\mem~31_combout ),
	.cout());
defparam \mem~31 .lut_mask = 16'hAACC;
defparam \mem~31 .sum_lutc_input = "datac";

dffeas \mem[5][2] (
	.clk(clk),
	.d(\mem~31_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\mem[5][2]~q ),
	.prn(vcc));
defparam \mem[5][2] .is_wysiwyg = "true";
defparam \mem[5][2] .power_up = "low";

cycloneive_lcell_comb \mem~25 (
	.dataa(\mem[5][2]~q ),
	.datab(src_channel_2),
	.datac(gnd),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\mem~25_combout ),
	.cout());
defparam \mem~25 .lut_mask = 16'hAACC;
defparam \mem~25 .sum_lutc_input = "datac";

dffeas \mem[4][2] (
	.clk(clk),
	.d(\mem~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(\mem[4][2]~q ),
	.prn(vcc));
defparam \mem[4][2] .is_wysiwyg = "true";
defparam \mem[4][2] .power_up = "low";

cycloneive_lcell_comb \mem~19 (
	.dataa(\mem[4][2]~q ),
	.datab(src_channel_2),
	.datac(gnd),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\mem~19_combout ),
	.cout());
defparam \mem~19 .lut_mask = 16'hAACC;
defparam \mem~19 .sum_lutc_input = "datac";

dffeas \mem[3][2] (
	.clk(clk),
	.d(\mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\mem[3][2]~q ),
	.prn(vcc));
defparam \mem[3][2] .is_wysiwyg = "true";
defparam \mem[3][2] .power_up = "low";

cycloneive_lcell_comb \mem~13 (
	.dataa(\mem[3][2]~q ),
	.datab(src_channel_2),
	.datac(gnd),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\mem~13_combout ),
	.cout());
defparam \mem~13 .lut_mask = 16'hAACC;
defparam \mem~13 .sum_lutc_input = "datac";

dffeas \mem[2][2] (
	.clk(clk),
	.d(\mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(\mem[2][2]~q ),
	.prn(vcc));
defparam \mem[2][2] .is_wysiwyg = "true";
defparam \mem[2][2] .power_up = "low";

cycloneive_lcell_comb \mem~7 (
	.dataa(\mem[2][2]~q ),
	.datab(src_channel_2),
	.datac(gnd),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\mem~7_combout ),
	.cout());
defparam \mem~7 .lut_mask = 16'hAACC;
defparam \mem~7 .sum_lutc_input = "datac";

dffeas \mem[1][2] (
	.clk(clk),
	.d(\mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\mem[1][2]~q ),
	.prn(vcc));
defparam \mem[1][2] .is_wysiwyg = "true";
defparam \mem[1][2] .power_up = "low";

cycloneive_lcell_comb \mem~1 (
	.dataa(\mem[1][2]~q ),
	.datab(src_channel_2),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~1_combout ),
	.cout());
defparam \mem~1 .lut_mask = 16'hAACC;
defparam \mem~1 .sum_lutc_input = "datac";

dffeas \mem[0][2] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\internal_out_valid~0_combout ),
	.q(\mem[0][2]~q ),
	.prn(vcc));
defparam \mem[0][2] .is_wysiwyg = "true";
defparam \mem[0][2] .power_up = "low";

dffeas \mem[9][1] (
	.clk(clk),
	.d(\mem~50_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[9][1]~q ),
	.prn(vcc));
defparam \mem[9][1] .is_wysiwyg = "true";
defparam \mem[9][1] .power_up = "low";

cycloneive_lcell_comb \mem~50 (
	.dataa(\mem[9][1]~q ),
	.datab(src_channel_1),
	.datac(gnd),
	.datad(mem_used_9),
	.cin(gnd),
	.combout(\mem~50_combout ),
	.cout());
defparam \mem~50 .lut_mask = 16'hAACC;
defparam \mem~50 .sum_lutc_input = "datac";

dffeas \mem[8][1] (
	.clk(clk),
	.d(\mem~50_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always8~0_combout ),
	.q(\mem[8][1]~q ),
	.prn(vcc));
defparam \mem[8][1] .is_wysiwyg = "true";
defparam \mem[8][1] .power_up = "low";

cycloneive_lcell_comb \mem~44 (
	.dataa(\mem[8][1]~q ),
	.datab(src_channel_1),
	.datac(gnd),
	.datad(\mem_used[8]~q ),
	.cin(gnd),
	.combout(\mem~44_combout ),
	.cout());
defparam \mem~44 .lut_mask = 16'hAACC;
defparam \mem~44 .sum_lutc_input = "datac";

dffeas \mem[7][1] (
	.clk(clk),
	.d(\mem~44_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\mem[7][1]~q ),
	.prn(vcc));
defparam \mem[7][1] .is_wysiwyg = "true";
defparam \mem[7][1] .power_up = "low";

cycloneive_lcell_comb \mem~38 (
	.dataa(\mem[7][1]~q ),
	.datab(src_channel_1),
	.datac(gnd),
	.datad(\mem_used[7]~q ),
	.cin(gnd),
	.combout(\mem~38_combout ),
	.cout());
defparam \mem~38 .lut_mask = 16'hAACC;
defparam \mem~38 .sum_lutc_input = "datac";

dffeas \mem[6][1] (
	.clk(clk),
	.d(\mem~38_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][1]~q ),
	.prn(vcc));
defparam \mem[6][1] .is_wysiwyg = "true";
defparam \mem[6][1] .power_up = "low";

cycloneive_lcell_comb \mem~32 (
	.dataa(\mem[6][1]~q ),
	.datab(src_channel_1),
	.datac(gnd),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\mem~32_combout ),
	.cout());
defparam \mem~32 .lut_mask = 16'hAACC;
defparam \mem~32 .sum_lutc_input = "datac";

dffeas \mem[5][1] (
	.clk(clk),
	.d(\mem~32_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\mem[5][1]~q ),
	.prn(vcc));
defparam \mem[5][1] .is_wysiwyg = "true";
defparam \mem[5][1] .power_up = "low";

cycloneive_lcell_comb \mem~26 (
	.dataa(\mem[5][1]~q ),
	.datab(src_channel_1),
	.datac(gnd),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\mem~26_combout ),
	.cout());
defparam \mem~26 .lut_mask = 16'hAACC;
defparam \mem~26 .sum_lutc_input = "datac";

dffeas \mem[4][1] (
	.clk(clk),
	.d(\mem~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(\mem[4][1]~q ),
	.prn(vcc));
defparam \mem[4][1] .is_wysiwyg = "true";
defparam \mem[4][1] .power_up = "low";

cycloneive_lcell_comb \mem~20 (
	.dataa(\mem[4][1]~q ),
	.datab(src_channel_1),
	.datac(gnd),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\mem~20_combout ),
	.cout());
defparam \mem~20 .lut_mask = 16'hAACC;
defparam \mem~20 .sum_lutc_input = "datac";

dffeas \mem[3][1] (
	.clk(clk),
	.d(\mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\mem[3][1]~q ),
	.prn(vcc));
defparam \mem[3][1] .is_wysiwyg = "true";
defparam \mem[3][1] .power_up = "low";

cycloneive_lcell_comb \mem~14 (
	.dataa(\mem[3][1]~q ),
	.datab(src_channel_1),
	.datac(gnd),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\mem~14_combout ),
	.cout());
defparam \mem~14 .lut_mask = 16'hAACC;
defparam \mem~14 .sum_lutc_input = "datac";

dffeas \mem[2][1] (
	.clk(clk),
	.d(\mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(\mem[2][1]~q ),
	.prn(vcc));
defparam \mem[2][1] .is_wysiwyg = "true";
defparam \mem[2][1] .power_up = "low";

cycloneive_lcell_comb \mem~8 (
	.dataa(\mem[2][1]~q ),
	.datab(src_channel_1),
	.datac(gnd),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\mem~8_combout ),
	.cout());
defparam \mem~8 .lut_mask = 16'hAACC;
defparam \mem~8 .sum_lutc_input = "datac";

dffeas \mem[1][1] (
	.clk(clk),
	.d(\mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\mem[1][1]~q ),
	.prn(vcc));
defparam \mem[1][1] .is_wysiwyg = "true";
defparam \mem[1][1] .power_up = "low";

cycloneive_lcell_comb \mem~2 (
	.dataa(\mem[1][1]~q ),
	.datab(src_channel_1),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'hAACC;
defparam \mem~2 .sum_lutc_input = "datac";

dffeas \mem[0][1] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\internal_out_valid~0_combout ),
	.q(\mem[0][1]~q ),
	.prn(vcc));
defparam \mem[0][1] .is_wysiwyg = "true";
defparam \mem[0][1] .power_up = "low";

dffeas \mem[9][0] (
	.clk(clk),
	.d(\mem~51_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[9][0]~q ),
	.prn(vcc));
defparam \mem[9][0] .is_wysiwyg = "true";
defparam \mem[9][0] .power_up = "low";

cycloneive_lcell_comb \mem~51 (
	.dataa(\mem[9][0]~q ),
	.datab(src_channel_0),
	.datac(gnd),
	.datad(mem_used_9),
	.cin(gnd),
	.combout(\mem~51_combout ),
	.cout());
defparam \mem~51 .lut_mask = 16'hAACC;
defparam \mem~51 .sum_lutc_input = "datac";

dffeas \mem[8][0] (
	.clk(clk),
	.d(\mem~51_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always8~0_combout ),
	.q(\mem[8][0]~q ),
	.prn(vcc));
defparam \mem[8][0] .is_wysiwyg = "true";
defparam \mem[8][0] .power_up = "low";

cycloneive_lcell_comb \mem~45 (
	.dataa(\mem[8][0]~q ),
	.datab(src_channel_0),
	.datac(gnd),
	.datad(\mem_used[8]~q ),
	.cin(gnd),
	.combout(\mem~45_combout ),
	.cout());
defparam \mem~45 .lut_mask = 16'hAACC;
defparam \mem~45 .sum_lutc_input = "datac";

dffeas \mem[7][0] (
	.clk(clk),
	.d(\mem~45_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\mem[7][0]~q ),
	.prn(vcc));
defparam \mem[7][0] .is_wysiwyg = "true";
defparam \mem[7][0] .power_up = "low";

cycloneive_lcell_comb \mem~39 (
	.dataa(\mem[7][0]~q ),
	.datab(src_channel_0),
	.datac(gnd),
	.datad(\mem_used[7]~q ),
	.cin(gnd),
	.combout(\mem~39_combout ),
	.cout());
defparam \mem~39 .lut_mask = 16'hAACC;
defparam \mem~39 .sum_lutc_input = "datac";

dffeas \mem[6][0] (
	.clk(clk),
	.d(\mem~39_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][0]~q ),
	.prn(vcc));
defparam \mem[6][0] .is_wysiwyg = "true";
defparam \mem[6][0] .power_up = "low";

cycloneive_lcell_comb \mem~33 (
	.dataa(\mem[6][0]~q ),
	.datab(src_channel_0),
	.datac(gnd),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\mem~33_combout ),
	.cout());
defparam \mem~33 .lut_mask = 16'hAACC;
defparam \mem~33 .sum_lutc_input = "datac";

dffeas \mem[5][0] (
	.clk(clk),
	.d(\mem~33_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\mem[5][0]~q ),
	.prn(vcc));
defparam \mem[5][0] .is_wysiwyg = "true";
defparam \mem[5][0] .power_up = "low";

cycloneive_lcell_comb \mem~27 (
	.dataa(\mem[5][0]~q ),
	.datab(src_channel_0),
	.datac(gnd),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\mem~27_combout ),
	.cout());
defparam \mem~27 .lut_mask = 16'hAACC;
defparam \mem~27 .sum_lutc_input = "datac";

dffeas \mem[4][0] (
	.clk(clk),
	.d(\mem~27_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(\mem[4][0]~q ),
	.prn(vcc));
defparam \mem[4][0] .is_wysiwyg = "true";
defparam \mem[4][0] .power_up = "low";

cycloneive_lcell_comb \mem~21 (
	.dataa(\mem[4][0]~q ),
	.datab(src_channel_0),
	.datac(gnd),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\mem~21_combout ),
	.cout());
defparam \mem~21 .lut_mask = 16'hAACC;
defparam \mem~21 .sum_lutc_input = "datac";

dffeas \mem[3][0] (
	.clk(clk),
	.d(\mem~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\mem[3][0]~q ),
	.prn(vcc));
defparam \mem[3][0] .is_wysiwyg = "true";
defparam \mem[3][0] .power_up = "low";

cycloneive_lcell_comb \mem~15 (
	.dataa(\mem[3][0]~q ),
	.datab(src_channel_0),
	.datac(gnd),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\mem~15_combout ),
	.cout());
defparam \mem~15 .lut_mask = 16'hAACC;
defparam \mem~15 .sum_lutc_input = "datac";

dffeas \mem[2][0] (
	.clk(clk),
	.d(\mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(\mem[2][0]~q ),
	.prn(vcc));
defparam \mem[2][0] .is_wysiwyg = "true";
defparam \mem[2][0] .power_up = "low";

cycloneive_lcell_comb \mem~9 (
	.dataa(\mem[2][0]~q ),
	.datab(src_channel_0),
	.datac(gnd),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\mem~9_combout ),
	.cout());
defparam \mem~9 .lut_mask = 16'hAACC;
defparam \mem~9 .sum_lutc_input = "datac";

dffeas \mem[1][0] (
	.clk(clk),
	.d(\mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\mem[1][0]~q ),
	.prn(vcc));
defparam \mem[1][0] .is_wysiwyg = "true";
defparam \mem[1][0] .power_up = "low";

cycloneive_lcell_comb \mem~3 (
	.dataa(\mem[1][0]~q ),
	.datab(src_channel_0),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~3_combout ),
	.cout());
defparam \mem~3 .lut_mask = 16'hAACC;
defparam \mem~3 .sum_lutc_input = "datac";

dffeas \mem[0][0] (
	.clk(clk),
	.d(\mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\internal_out_valid~0_combout ),
	.q(\mem[0][0]~q ),
	.prn(vcc));
defparam \mem[0][0] .is_wysiwyg = "true";
defparam \mem[0][0] .power_up = "low";

cycloneive_lcell_comb \mem_used[9]~0 (
	.dataa(\read~0_combout ),
	.datab(mem_used_9),
	.datac(WideOr1),
	.datad(\mem_used[8]~q ),
	.cin(gnd),
	.combout(\mem_used[9]~0_combout ),
	.cout());
defparam \mem_used[9]~0 .lut_mask = 16'hA888;
defparam \mem_used[9]~0 .sum_lutc_input = "datac";

dffeas \mem[9][16] (
	.clk(clk),
	.d(\mem~52_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[9][16]~q ),
	.prn(vcc));
defparam \mem[9][16] .is_wysiwyg = "true";
defparam \mem[9][16] .power_up = "low";

cycloneive_lcell_comb \mem~52 (
	.dataa(\mem[9][16]~q ),
	.datab(src_payload_0),
	.datac(gnd),
	.datad(mem_used_9),
	.cin(gnd),
	.combout(\mem~52_combout ),
	.cout());
defparam \mem~52 .lut_mask = 16'hAACC;
defparam \mem~52 .sum_lutc_input = "datac";

dffeas \mem[8][16] (
	.clk(clk),
	.d(\mem~52_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always8~0_combout ),
	.q(\mem[8][16]~q ),
	.prn(vcc));
defparam \mem[8][16] .is_wysiwyg = "true";
defparam \mem[8][16] .power_up = "low";

cycloneive_lcell_comb \mem~46 (
	.dataa(\mem[8][16]~q ),
	.datab(src_payload_0),
	.datac(gnd),
	.datad(\mem_used[8]~q ),
	.cin(gnd),
	.combout(\mem~46_combout ),
	.cout());
defparam \mem~46 .lut_mask = 16'hAACC;
defparam \mem~46 .sum_lutc_input = "datac";

dffeas \mem[7][16] (
	.clk(clk),
	.d(\mem~46_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\mem[7][16]~q ),
	.prn(vcc));
defparam \mem[7][16] .is_wysiwyg = "true";
defparam \mem[7][16] .power_up = "low";

cycloneive_lcell_comb \mem~40 (
	.dataa(\mem[7][16]~q ),
	.datab(src_payload_0),
	.datac(gnd),
	.datad(\mem_used[7]~q ),
	.cin(gnd),
	.combout(\mem~40_combout ),
	.cout());
defparam \mem~40 .lut_mask = 16'hAACC;
defparam \mem~40 .sum_lutc_input = "datac";

dffeas \mem[6][16] (
	.clk(clk),
	.d(\mem~40_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][16]~q ),
	.prn(vcc));
defparam \mem[6][16] .is_wysiwyg = "true";
defparam \mem[6][16] .power_up = "low";

cycloneive_lcell_comb \mem~34 (
	.dataa(\mem[6][16]~q ),
	.datab(src_payload_0),
	.datac(gnd),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\mem~34_combout ),
	.cout());
defparam \mem~34 .lut_mask = 16'hAACC;
defparam \mem~34 .sum_lutc_input = "datac";

dffeas \mem[5][16] (
	.clk(clk),
	.d(\mem~34_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\mem[5][16]~q ),
	.prn(vcc));
defparam \mem[5][16] .is_wysiwyg = "true";
defparam \mem[5][16] .power_up = "low";

cycloneive_lcell_comb \mem~28 (
	.dataa(\mem[5][16]~q ),
	.datab(src_payload_0),
	.datac(gnd),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\mem~28_combout ),
	.cout());
defparam \mem~28 .lut_mask = 16'hAACC;
defparam \mem~28 .sum_lutc_input = "datac";

dffeas \mem[4][16] (
	.clk(clk),
	.d(\mem~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(\mem[4][16]~q ),
	.prn(vcc));
defparam \mem[4][16] .is_wysiwyg = "true";
defparam \mem[4][16] .power_up = "low";

cycloneive_lcell_comb \mem~22 (
	.dataa(\mem[4][16]~q ),
	.datab(src_payload_0),
	.datac(gnd),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\mem~22_combout ),
	.cout());
defparam \mem~22 .lut_mask = 16'hAACC;
defparam \mem~22 .sum_lutc_input = "datac";

dffeas \mem[3][16] (
	.clk(clk),
	.d(\mem~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\mem[3][16]~q ),
	.prn(vcc));
defparam \mem[3][16] .is_wysiwyg = "true";
defparam \mem[3][16] .power_up = "low";

cycloneive_lcell_comb \mem~16 (
	.dataa(\mem[3][16]~q ),
	.datab(src_payload_0),
	.datac(gnd),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\mem~16_combout ),
	.cout());
defparam \mem~16 .lut_mask = 16'hAACC;
defparam \mem~16 .sum_lutc_input = "datac";

dffeas \mem[2][16] (
	.clk(clk),
	.d(\mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(\mem[2][16]~q ),
	.prn(vcc));
defparam \mem[2][16] .is_wysiwyg = "true";
defparam \mem[2][16] .power_up = "low";

cycloneive_lcell_comb \mem~10 (
	.dataa(\mem[2][16]~q ),
	.datab(src_payload_0),
	.datac(gnd),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\mem~10_combout ),
	.cout());
defparam \mem~10 .lut_mask = 16'hAACC;
defparam \mem~10 .sum_lutc_input = "datac";

dffeas \mem[1][16] (
	.clk(clk),
	.d(\mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\mem[1][16]~q ),
	.prn(vcc));
defparam \mem[1][16] .is_wysiwyg = "true";
defparam \mem[1][16] .power_up = "low";

cycloneive_lcell_comb \mem~4 (
	.dataa(\mem[1][16]~q ),
	.datab(src_payload_0),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~4_combout ),
	.cout());
defparam \mem~4 .lut_mask = 16'hAACC;
defparam \mem~4 .sum_lutc_input = "datac";

dffeas \mem[0][16] (
	.clk(clk),
	.d(\mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\internal_out_valid~0_combout ),
	.q(\mem[0][16]~q ),
	.prn(vcc));
defparam \mem[0][16] .is_wysiwyg = "true";
defparam \mem[0][16] .power_up = "low";

dffeas \mem[9][8] (
	.clk(clk),
	.d(\mem~53_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[9][8]~q ),
	.prn(vcc));
defparam \mem[9][8] .is_wysiwyg = "true";
defparam \mem[9][8] .power_up = "low";

cycloneive_lcell_comb \mem~53 (
	.dataa(\mem[9][8]~q ),
	.datab(src_channel_8),
	.datac(gnd),
	.datad(mem_used_9),
	.cin(gnd),
	.combout(\mem~53_combout ),
	.cout());
defparam \mem~53 .lut_mask = 16'hAACC;
defparam \mem~53 .sum_lutc_input = "datac";

dffeas \mem[8][8] (
	.clk(clk),
	.d(\mem~53_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always8~0_combout ),
	.q(\mem[8][8]~q ),
	.prn(vcc));
defparam \mem[8][8] .is_wysiwyg = "true";
defparam \mem[8][8] .power_up = "low";

cycloneive_lcell_comb \mem~47 (
	.dataa(\mem[8][8]~q ),
	.datab(src_channel_8),
	.datac(gnd),
	.datad(\mem_used[8]~q ),
	.cin(gnd),
	.combout(\mem~47_combout ),
	.cout());
defparam \mem~47 .lut_mask = 16'hAACC;
defparam \mem~47 .sum_lutc_input = "datac";

dffeas \mem[7][8] (
	.clk(clk),
	.d(\mem~47_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always7~0_combout ),
	.q(\mem[7][8]~q ),
	.prn(vcc));
defparam \mem[7][8] .is_wysiwyg = "true";
defparam \mem[7][8] .power_up = "low";

cycloneive_lcell_comb \mem~41 (
	.dataa(\mem[7][8]~q ),
	.datab(src_channel_8),
	.datac(gnd),
	.datad(\mem_used[7]~q ),
	.cin(gnd),
	.combout(\mem~41_combout ),
	.cout());
defparam \mem~41 .lut_mask = 16'hAACC;
defparam \mem~41 .sum_lutc_input = "datac";

dffeas \mem[6][8] (
	.clk(clk),
	.d(\mem~41_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always6~0_combout ),
	.q(\mem[6][8]~q ),
	.prn(vcc));
defparam \mem[6][8] .is_wysiwyg = "true";
defparam \mem[6][8] .power_up = "low";

cycloneive_lcell_comb \mem~35 (
	.dataa(\mem[6][8]~q ),
	.datab(src_channel_8),
	.datac(gnd),
	.datad(\mem_used[6]~q ),
	.cin(gnd),
	.combout(\mem~35_combout ),
	.cout());
defparam \mem~35 .lut_mask = 16'hAACC;
defparam \mem~35 .sum_lutc_input = "datac";

dffeas \mem[5][8] (
	.clk(clk),
	.d(\mem~35_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always5~0_combout ),
	.q(\mem[5][8]~q ),
	.prn(vcc));
defparam \mem[5][8] .is_wysiwyg = "true";
defparam \mem[5][8] .power_up = "low";

cycloneive_lcell_comb \mem~29 (
	.dataa(\mem[5][8]~q ),
	.datab(src_channel_8),
	.datac(gnd),
	.datad(\mem_used[5]~q ),
	.cin(gnd),
	.combout(\mem~29_combout ),
	.cout());
defparam \mem~29 .lut_mask = 16'hAACC;
defparam \mem~29 .sum_lutc_input = "datac";

dffeas \mem[4][8] (
	.clk(clk),
	.d(\mem~29_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(\mem[4][8]~q ),
	.prn(vcc));
defparam \mem[4][8] .is_wysiwyg = "true";
defparam \mem[4][8] .power_up = "low";

cycloneive_lcell_comb \mem~23 (
	.dataa(\mem[4][8]~q ),
	.datab(src_channel_8),
	.datac(gnd),
	.datad(\mem_used[4]~q ),
	.cin(gnd),
	.combout(\mem~23_combout ),
	.cout());
defparam \mem~23 .lut_mask = 16'hAACC;
defparam \mem~23 .sum_lutc_input = "datac";

dffeas \mem[3][8] (
	.clk(clk),
	.d(\mem~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\mem[3][8]~q ),
	.prn(vcc));
defparam \mem[3][8] .is_wysiwyg = "true";
defparam \mem[3][8] .power_up = "low";

cycloneive_lcell_comb \mem~17 (
	.dataa(\mem[3][8]~q ),
	.datab(src_channel_8),
	.datac(gnd),
	.datad(\mem_used[3]~q ),
	.cin(gnd),
	.combout(\mem~17_combout ),
	.cout());
defparam \mem~17 .lut_mask = 16'hAACC;
defparam \mem~17 .sum_lutc_input = "datac";

dffeas \mem[2][8] (
	.clk(clk),
	.d(\mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always2~0_combout ),
	.q(\mem[2][8]~q ),
	.prn(vcc));
defparam \mem[2][8] .is_wysiwyg = "true";
defparam \mem[2][8] .power_up = "low";

cycloneive_lcell_comb \mem~11 (
	.dataa(\mem[2][8]~q ),
	.datab(src_channel_8),
	.datac(gnd),
	.datad(\mem_used[2]~q ),
	.cin(gnd),
	.combout(\mem~11_combout ),
	.cout());
defparam \mem~11 .lut_mask = 16'hAACC;
defparam \mem~11 .sum_lutc_input = "datac";

dffeas \mem[1][8] (
	.clk(clk),
	.d(\mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\mem[1][8]~q ),
	.prn(vcc));
defparam \mem[1][8] .is_wysiwyg = "true";
defparam \mem[1][8] .power_up = "low";

cycloneive_lcell_comb \mem~5 (
	.dataa(\mem[1][8]~q ),
	.datab(src_channel_8),
	.datac(gnd),
	.datad(\mem_used[1]~q ),
	.cin(gnd),
	.combout(\mem~5_combout ),
	.cout());
defparam \mem~5 .lut_mask = 16'hAACC;
defparam \mem~5 .sum_lutc_input = "datac";

dffeas \mem[0][8] (
	.clk(clk),
	.d(\mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\internal_out_valid~0_combout ),
	.q(\mem[0][8]~q ),
	.prn(vcc));
defparam \mem[0][8] .is_wysiwyg = "true";
defparam \mem[0][8] .power_up = "low";

endmodule

module flashLoader_qspi_inf_mux (
	altera_reset_synchronizer_int_chain_out,
	out_valid,
	grant_0,
	out_valid1,
	out_valid2,
	request_1,
	full_addercout_1,
	cout,
	sum_1,
	request_2,
	cout1,
	grant_01,
	WideOr1,
	write,
	out_endofpacket,
	out_endofpacket1,
	out_endofpacket2,
	src_payload_0,
	out_data_0,
	out_data_01,
	out_data_02,
	src_data_0,
	out_channel_2,
	out_channel_21,
	out_channel_22,
	src_channel_2,
	out_channel_1,
	out_channel_11,
	out_channel_12,
	src_channel_1,
	out_channel_0,
	out_channel_01,
	out_channel_02,
	src_channel_0,
	out_channel_8,
	out_channel_81,
	out_channel_82,
	src_channel_8,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	altera_reset_synchronizer_int_chain_out;
input 	out_valid;
output 	grant_0;
input 	out_valid1;
input 	out_valid2;
output 	request_1;
output 	full_addercout_1;
output 	cout;
output 	sum_1;
output 	request_2;
output 	cout1;
output 	grant_01;
output 	WideOr1;
input 	write;
input 	out_endofpacket;
input 	out_endofpacket1;
input 	out_endofpacket2;
output 	src_payload_0;
input 	out_data_0;
input 	out_data_01;
input 	out_data_02;
output 	src_data_0;
input 	out_channel_2;
input 	out_channel_21;
input 	out_channel_22;
output 	src_channel_2;
input 	out_channel_1;
input 	out_channel_11;
input 	out_channel_12;
output 	src_channel_1;
input 	out_channel_0;
input 	out_channel_01;
input 	out_channel_02;
output 	src_channel_0;
input 	out_channel_8;
input 	out_channel_81;
input 	out_channel_82;
output 	src_channel_8;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



flashLoader_flashLoader_intel_generic_serial_flash_interface_top_0_qspi_inf_inst_qspi_inf_mux_qspi_inf_mux qspi_inf_mux(
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.out_valid(out_valid),
	.grant_0(grant_0),
	.out_valid1(out_valid1),
	.out_valid2(out_valid2),
	.request_1(request_1),
	.full_addercout_1(full_addercout_1),
	.cout(cout),
	.sum_1(sum_1),
	.request_2(request_2),
	.cout1(cout1),
	.grant_01(grant_01),
	.WideOr1(WideOr1),
	.write(write),
	.out_endofpacket(out_endofpacket),
	.out_endofpacket1(out_endofpacket1),
	.out_endofpacket2(out_endofpacket2),
	.src_payload_0(src_payload_0),
	.out_data_0(out_data_0),
	.out_data_01(out_data_01),
	.out_data_02(out_data_02),
	.src_data_0(src_data_0),
	.out_channel_2(out_channel_2),
	.out_channel_21(out_channel_21),
	.out_channel_22(out_channel_22),
	.src_channel_2(src_channel_2),
	.out_channel_1(out_channel_1),
	.out_channel_11(out_channel_11),
	.out_channel_12(out_channel_12),
	.src_channel_1(src_channel_1),
	.out_channel_0(out_channel_0),
	.out_channel_01(out_channel_01),
	.out_channel_02(out_channel_02),
	.src_channel_0(src_channel_0),
	.out_channel_8(out_channel_8),
	.out_channel_81(out_channel_81),
	.out_channel_82(out_channel_82),
	.src_channel_8(src_channel_8),
	.clk_clk(clk_clk));

endmodule

module flashLoader_flashLoader_intel_generic_serial_flash_interface_top_0_qspi_inf_inst_qspi_inf_mux_qspi_inf_mux (
	altera_reset_synchronizer_int_chain_out,
	out_valid,
	grant_0,
	out_valid1,
	out_valid2,
	request_1,
	full_addercout_1,
	cout,
	sum_1,
	request_2,
	cout1,
	grant_01,
	WideOr1,
	write,
	out_endofpacket,
	out_endofpacket1,
	out_endofpacket2,
	src_payload_0,
	out_data_0,
	out_data_01,
	out_data_02,
	src_data_0,
	out_channel_2,
	out_channel_21,
	out_channel_22,
	src_channel_2,
	out_channel_1,
	out_channel_11,
	out_channel_12,
	src_channel_1,
	out_channel_0,
	out_channel_01,
	out_channel_02,
	src_channel_0,
	out_channel_8,
	out_channel_81,
	out_channel_82,
	src_channel_8,
	clk_clk)/* synthesis synthesis_greybox=0 */;
input 	altera_reset_synchronizer_int_chain_out;
input 	out_valid;
output 	grant_0;
input 	out_valid1;
input 	out_valid2;
output 	request_1;
output 	full_addercout_1;
output 	cout;
output 	sum_1;
output 	request_2;
output 	cout1;
output 	grant_01;
output 	WideOr1;
input 	write;
input 	out_endofpacket;
input 	out_endofpacket1;
input 	out_endofpacket2;
output 	src_payload_0;
input 	out_data_0;
input 	out_data_01;
input 	out_data_02;
output 	src_data_0;
input 	out_channel_2;
input 	out_channel_21;
input 	out_channel_22;
output 	src_channel_2;
input 	out_channel_1;
input 	out_channel_11;
input 	out_channel_12;
output 	src_channel_1;
input 	out_channel_0;
input 	out_channel_01;
input 	out_channel_02;
output 	src_channel_0;
input 	out_channel_8;
input 	out_channel_81;
input 	out_channel_82;
output 	src_channel_8;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \prev_request[0]~q ;
wire \arb|grant[2]~4_combout ;
wire \arb|grant[2]~5_combout ;
wire \arb|grant[0]~6_combout ;
wire \prev_request[0]~1_combout ;
wire \arb|grant[1]~7_combout ;
wire \prev_request[1]~2_combout ;
wire \prev_request[1]~q ;
wire \prev_request[2]~0_combout ;
wire \prev_request[2]~q ;
wire \src_valid~0_combout ;
wire \WideOr1~3_combout ;
wire \src_payload[0]~0_combout ;
wire \src_data[0]~0_combout ;
wire \src_channel[2]~0_combout ;
wire \src_channel[1]~2_combout ;
wire \src_channel[0]~4_combout ;
wire \src_channel[8]~6_combout ;


flashLoader_altera_merlin_arbitrator_1 arb(
	.reset(altera_reset_synchronizer_int_chain_out),
	.out_valid(out_valid),
	.prev_request_2(\prev_request[2]~q ),
	.grant_0(grant_0),
	.out_valid1(out_valid1),
	.prev_request_0(\prev_request[0]~q ),
	.out_valid2(out_valid2),
	.prev_request_1(\prev_request[1]~q ),
	.request_1(request_1),
	.full_addercout_1(full_addercout_1),
	.cout(cout),
	.sum_1(sum_1),
	.request_2(request_2),
	.cout1(cout1),
	.grant_01(grant_01),
	.grant_2(\arb|grant[2]~4_combout ),
	.grant_21(\arb|grant[2]~5_combout ),
	.WideOr1(WideOr1),
	.write(write),
	.grant_02(\arb|grant[0]~6_combout ),
	.src_payload_0(src_payload_0),
	.grant_1(\arb|grant[1]~7_combout ),
	.clk(clk_clk));

dffeas \prev_request[0] (
	.clk(clk_clk),
	.d(\prev_request[0]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\prev_request[0]~q ),
	.prn(vcc));
defparam \prev_request[0] .is_wysiwyg = "true";
defparam \prev_request[0] .power_up = "low";

cycloneive_lcell_comb \prev_request[0]~1 (
	.dataa(\prev_request[0]~q ),
	.datab(gnd),
	.datac(out_valid1),
	.datad(out_endofpacket1),
	.cin(gnd),
	.combout(\prev_request[0]~1_combout ),
	.cout());
defparam \prev_request[0]~1 .lut_mask = 16'h0AFA;
defparam \prev_request[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \request[1] (
	.dataa(out_valid2),
	.datab(\prev_request[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(request_1),
	.cout());
defparam \request[1] .lut_mask = 16'hEEEE;
defparam \request[1] .sum_lutc_input = "datac";

cycloneive_lcell_comb \request[2] (
	.dataa(out_valid),
	.datab(\prev_request[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(request_2),
	.cout());
defparam \request[2] .lut_mask = 16'hEEEE;
defparam \request[2] .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr1~2 (
	.dataa(\src_valid~0_combout ),
	.datab(\WideOr1~3_combout ),
	.datac(out_valid),
	.datad(\arb|grant[2]~5_combout ),
	.cin(gnd),
	.combout(WideOr1),
	.cout());
defparam \WideOr1~2 .lut_mask = 16'hFEEE;
defparam \WideOr1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload[0]~1 (
	.dataa(\src_payload[0]~0_combout ),
	.datab(out_endofpacket2),
	.datac(\arb|grant[1]~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload_0),
	.cout());
defparam \src_payload[0]~1 .lut_mask = 16'hEAEA;
defparam \src_payload[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0]~1 (
	.dataa(\src_data[0]~0_combout ),
	.datab(\arb|grant[1]~7_combout ),
	.datac(out_data_02),
	.datad(gnd),
	.cin(gnd),
	.combout(src_data_0),
	.cout());
defparam \src_data[0]~1 .lut_mask = 16'hEAEA;
defparam \src_data[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[2]~1 (
	.dataa(\src_channel[2]~0_combout ),
	.datab(\arb|grant[1]~7_combout ),
	.datac(out_channel_22),
	.datad(gnd),
	.cin(gnd),
	.combout(src_channel_2),
	.cout());
defparam \src_channel[2]~1 .lut_mask = 16'hEAEA;
defparam \src_channel[2]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[1]~3 (
	.dataa(\src_channel[1]~2_combout ),
	.datab(\arb|grant[1]~7_combout ),
	.datac(out_channel_12),
	.datad(gnd),
	.cin(gnd),
	.combout(src_channel_1),
	.cout());
defparam \src_channel[1]~3 .lut_mask = 16'hEAEA;
defparam \src_channel[1]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[0]~5 (
	.dataa(\src_channel[0]~4_combout ),
	.datab(\arb|grant[1]~7_combout ),
	.datac(out_channel_02),
	.datad(gnd),
	.cin(gnd),
	.combout(src_channel_0),
	.cout());
defparam \src_channel[0]~5 .lut_mask = 16'hEAEA;
defparam \src_channel[0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[8]~7 (
	.dataa(\src_channel[8]~6_combout ),
	.datab(\arb|grant[1]~7_combout ),
	.datac(out_channel_82),
	.datad(gnd),
	.cin(gnd),
	.combout(src_channel_8),
	.cout());
defparam \src_channel[8]~7 .lut_mask = 16'hEAEA;
defparam \src_channel[8]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \prev_request[1]~2 (
	.dataa(\prev_request[1]~q ),
	.datab(gnd),
	.datac(out_valid2),
	.datad(out_endofpacket2),
	.cin(gnd),
	.combout(\prev_request[1]~2_combout ),
	.cout());
defparam \prev_request[1]~2 .lut_mask = 16'h0AFA;
defparam \prev_request[1]~2 .sum_lutc_input = "datac";

dffeas \prev_request[1] (
	.clk(clk_clk),
	.d(\prev_request[1]~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\prev_request[1]~q ),
	.prn(vcc));
defparam \prev_request[1] .is_wysiwyg = "true";
defparam \prev_request[1] .power_up = "low";

cycloneive_lcell_comb \prev_request[2]~0 (
	.dataa(\prev_request[2]~q ),
	.datab(gnd),
	.datac(out_valid),
	.datad(out_endofpacket),
	.cin(gnd),
	.combout(\prev_request[2]~0_combout ),
	.cout());
defparam \prev_request[2]~0 .lut_mask = 16'h0AFA;
defparam \prev_request[2]~0 .sum_lutc_input = "datac";

dffeas \prev_request[2] (
	.clk(clk_clk),
	.d(\prev_request[2]~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\prev_request[2]~q ),
	.prn(vcc));
defparam \prev_request[2] .is_wysiwyg = "true";
defparam \prev_request[2] .power_up = "low";

cycloneive_lcell_comb \src_valid~0 (
	.dataa(out_valid1),
	.datab(grant_0),
	.datac(full_addercout_1),
	.datad(cout),
	.cin(gnd),
	.combout(\src_valid~0_combout ),
	.cout());
defparam \src_valid~0 .lut_mask = 16'h88A8;
defparam \src_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \WideOr1~3 (
	.dataa(out_valid2),
	.datab(gnd),
	.datac(cout1),
	.datad(sum_1),
	.cin(gnd),
	.combout(\WideOr1~3_combout ),
	.cout());
defparam \WideOr1~3 .lut_mask = 16'hA0AA;
defparam \WideOr1~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_payload[0]~0 (
	.dataa(out_endofpacket),
	.datab(out_endofpacket1),
	.datac(\arb|grant[0]~6_combout ),
	.datad(\arb|grant[2]~4_combout ),
	.cin(gnd),
	.combout(\src_payload[0]~0_combout ),
	.cout());
defparam \src_payload[0]~0 .lut_mask = 16'hEAC0;
defparam \src_payload[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_data[0]~0 (
	.dataa(\arb|grant[0]~6_combout ),
	.datab(\arb|grant[2]~4_combout ),
	.datac(out_data_0),
	.datad(out_data_01),
	.cin(gnd),
	.combout(\src_data[0]~0_combout ),
	.cout());
defparam \src_data[0]~0 .lut_mask = 16'hEAC0;
defparam \src_data[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[2]~0 (
	.dataa(\arb|grant[0]~6_combout ),
	.datab(\arb|grant[2]~4_combout ),
	.datac(out_channel_2),
	.datad(out_channel_21),
	.cin(gnd),
	.combout(\src_channel[2]~0_combout ),
	.cout());
defparam \src_channel[2]~0 .lut_mask = 16'hEAC0;
defparam \src_channel[2]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[1]~2 (
	.dataa(\arb|grant[0]~6_combout ),
	.datab(\arb|grant[2]~4_combout ),
	.datac(out_channel_1),
	.datad(out_channel_11),
	.cin(gnd),
	.combout(\src_channel[1]~2_combout ),
	.cout());
defparam \src_channel[1]~2 .lut_mask = 16'hEAC0;
defparam \src_channel[1]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[0]~4 (
	.dataa(\arb|grant[0]~6_combout ),
	.datab(\arb|grant[2]~4_combout ),
	.datac(out_channel_0),
	.datad(out_channel_01),
	.cin(gnd),
	.combout(\src_channel[0]~4_combout ),
	.cout());
defparam \src_channel[0]~4 .lut_mask = 16'hEAC0;
defparam \src_channel[0]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \src_channel[8]~6 (
	.dataa(\arb|grant[0]~6_combout ),
	.datab(\arb|grant[2]~4_combout ),
	.datac(out_channel_8),
	.datad(out_channel_81),
	.cin(gnd),
	.combout(\src_channel[8]~6_combout ),
	.cout());
defparam \src_channel[8]~6 .lut_mask = 16'hEAC0;
defparam \src_channel[8]~6 .sum_lutc_input = "datac";

endmodule

module flashLoader_altera_merlin_arbitrator_1 (
	reset,
	out_valid,
	prev_request_2,
	grant_0,
	out_valid1,
	prev_request_0,
	out_valid2,
	prev_request_1,
	request_1,
	full_addercout_1,
	cout,
	sum_1,
	request_2,
	cout1,
	grant_01,
	grant_2,
	grant_21,
	WideOr1,
	write,
	grant_02,
	src_payload_0,
	grant_1,
	clk)/* synthesis synthesis_greybox=0 */;
input 	reset;
input 	out_valid;
input 	prev_request_2;
output 	grant_0;
input 	out_valid1;
input 	prev_request_0;
input 	out_valid2;
input 	prev_request_1;
input 	request_1;
output 	full_addercout_1;
output 	cout;
output 	sum_1;
input 	request_2;
output 	cout1;
output 	grant_01;
output 	grant_2;
output 	grant_21;
input 	WideOr1;
input 	write;
output 	grant_02;
input 	src_payload_0;
output 	grant_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \adder|full_adder.cout[0]~0_combout ;
wire \adder|sum[2]~combout ;
wire \WideOr0~combout ;
wire \top_priority_reg~2_combout ;
wire \top_priority_reg~3_combout ;
wire \top_priority_reg~4_combout ;
wire \top_priority_reg[0]~q ;
wire \top_priority_reg~5_combout ;
wire \top_priority_reg~6_combout ;
wire \top_priority_reg[1]~q ;
wire \top_priority_reg~0_combout ;
wire \top_priority_reg~1_combout ;
wire \top_priority_reg[2]~q ;


flashLoader_altera_merlin_arb_adder_1 adder(
	.top_priority_reg_2(\top_priority_reg[2]~q ),
	.out_valid(out_valid),
	.prev_request_2(prev_request_2),
	.top_priority_reg_0(\top_priority_reg[0]~q ),
	.top_priority_reg_1(\top_priority_reg[1]~q ),
	.out_valid1(out_valid1),
	.prev_request_0(prev_request_0),
	.full_addercout_0(\adder|full_adder.cout[0]~0_combout ),
	.request_1(request_1),
	.full_addercout_1(full_addercout_1),
	.cout(cout),
	.sum_1(sum_1),
	.request_2(request_2),
	.cout1(cout1),
	.sum_2(\adder|sum[2]~combout ));

cycloneive_lcell_comb \grant[0]~2 (
	.dataa(\top_priority_reg[2]~q ),
	.datab(out_valid),
	.datac(prev_request_2),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_0),
	.cout());
defparam \grant[0]~2 .lut_mask = 16'h02FF;
defparam \grant[0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \grant[0]~3 (
	.dataa(\top_priority_reg[2]~q ),
	.datab(full_addercout_1),
	.datac(request_2),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(grant_01),
	.cout());
defparam \grant[0]~3 .lut_mask = 16'h8EFF;
defparam \grant[0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \grant[2]~4 (
	.dataa(request_2),
	.datab(cout1),
	.datac(request_1),
	.datad(\adder|sum[2]~combout ),
	.cin(gnd),
	.combout(grant_2),
	.cout());
defparam \grant[2]~4 .lut_mask = 16'h08AA;
defparam \grant[2]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \grant[2]~5 (
	.dataa(cout1),
	.datab(request_1),
	.datac(request_2),
	.datad(\adder|sum[2]~combout ),
	.cin(gnd),
	.combout(grant_21),
	.cout());
defparam \grant[2]~5 .lut_mask = 16'h2DFF;
defparam \grant[2]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \grant[0]~6 (
	.dataa(grant_0),
	.datab(full_addercout_1),
	.datac(cout),
	.datad(\adder|full_adder.cout[0]~0_combout ),
	.cin(gnd),
	.combout(grant_02),
	.cout());
defparam \grant[0]~6 .lut_mask = 16'h00AE;
defparam \grant[0]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \grant[1]~7 (
	.dataa(out_valid2),
	.datab(prev_request_1),
	.datac(cout1),
	.datad(sum_1),
	.cin(gnd),
	.combout(grant_1),
	.cout());
defparam \grant[1]~7 .lut_mask = 16'hE0EE;
defparam \grant[1]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb WideOr0(
	.dataa(out_valid),
	.datab(prev_request_2),
	.datac(request_1),
	.datad(\adder|full_adder.cout[0]~0_combout ),
	.cin(gnd),
	.combout(\WideOr0~combout ),
	.cout());
defparam WideOr0.lut_mask = 16'hFEFF;
defparam WideOr0.sum_lutc_input = "datac";

cycloneive_lcell_comb \top_priority_reg~2 (
	.dataa(grant_2),
	.datab(\top_priority_reg[2]~q ),
	.datac(gnd),
	.datad(\WideOr0~combout ),
	.cin(gnd),
	.combout(\top_priority_reg~2_combout ),
	.cout());
defparam \top_priority_reg~2 .lut_mask = 16'hAACC;
defparam \top_priority_reg~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \top_priority_reg~3 (
	.dataa(grant_02),
	.datab(WideOr1),
	.datac(gnd),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(\top_priority_reg~3_combout ),
	.cout());
defparam \top_priority_reg~3 .lut_mask = 16'h88BB;
defparam \top_priority_reg~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \top_priority_reg~4 (
	.dataa(\top_priority_reg~2_combout ),
	.datab(\top_priority_reg~3_combout ),
	.datac(write),
	.datad(src_payload_0),
	.cin(gnd),
	.combout(\top_priority_reg~4_combout ),
	.cout());
defparam \top_priority_reg~4 .lut_mask = 16'h5333;
defparam \top_priority_reg~4 .sum_lutc_input = "datac";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

cycloneive_lcell_comb \top_priority_reg~5 (
	.dataa(grant_02),
	.datab(\WideOr0~combout ),
	.datac(gnd),
	.datad(\top_priority_reg[0]~q ),
	.cin(gnd),
	.combout(\top_priority_reg~5_combout ),
	.cout());
defparam \top_priority_reg~5 .lut_mask = 16'h88BB;
defparam \top_priority_reg~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \top_priority_reg~6 (
	.dataa(\top_priority_reg~5_combout ),
	.datab(grant_1),
	.datac(write),
	.datad(src_payload_0),
	.cin(gnd),
	.combout(\top_priority_reg~6_combout ),
	.cout());
defparam \top_priority_reg~6 .lut_mask = 16'hACCC;
defparam \top_priority_reg~6 .sum_lutc_input = "datac";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(\top_priority_reg~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(WideOr1),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

cycloneive_lcell_comb \top_priority_reg~0 (
	.dataa(grant_1),
	.datab(\top_priority_reg[1]~q ),
	.datac(gnd),
	.datad(\WideOr0~combout ),
	.cin(gnd),
	.combout(\top_priority_reg~0_combout ),
	.cout());
defparam \top_priority_reg~0 .lut_mask = 16'hAACC;
defparam \top_priority_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \top_priority_reg~1 (
	.dataa(\top_priority_reg~0_combout ),
	.datab(grant_2),
	.datac(write),
	.datad(src_payload_0),
	.cin(gnd),
	.combout(\top_priority_reg~1_combout ),
	.cout());
defparam \top_priority_reg~1 .lut_mask = 16'hACCC;
defparam \top_priority_reg~1 .sum_lutc_input = "datac";

dffeas \top_priority_reg[2] (
	.clk(clk),
	.d(\top_priority_reg~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(WideOr1),
	.q(\top_priority_reg[2]~q ),
	.prn(vcc));
defparam \top_priority_reg[2] .is_wysiwyg = "true";
defparam \top_priority_reg[2] .power_up = "low";

endmodule

module flashLoader_altera_merlin_arb_adder_1 (
	top_priority_reg_2,
	out_valid,
	prev_request_2,
	top_priority_reg_0,
	top_priority_reg_1,
	out_valid1,
	prev_request_0,
	full_addercout_0,
	request_1,
	full_addercout_1,
	cout,
	sum_1,
	request_2,
	cout1,
	sum_2)/* synthesis synthesis_greybox=0 */;
input 	top_priority_reg_2;
input 	out_valid;
input 	prev_request_2;
input 	top_priority_reg_0;
input 	top_priority_reg_1;
input 	out_valid1;
input 	prev_request_0;
output 	full_addercout_0;
input 	request_1;
output 	full_addercout_1;
output 	cout;
output 	sum_1;
input 	request_2;
output 	cout1;
output 	sum_2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneive_lcell_comb \full_adder.cout[0]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(out_valid1),
	.datad(prev_request_0),
	.cin(gnd),
	.combout(full_addercout_0),
	.cout());
defparam \full_adder.cout[0]~0 .lut_mask = 16'h000F;
defparam \full_adder.cout[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \full_adder.cout[1] (
	.dataa(top_priority_reg_1),
	.datab(full_addercout_0),
	.datac(top_priority_reg_0),
	.datad(request_1),
	.cin(gnd),
	.combout(full_addercout_1),
	.cout());
defparam \full_adder.cout[1] .lut_mask = 16'h08AE;
defparam \full_adder.cout[1] .sum_lutc_input = "datac";

cycloneive_lcell_comb \cout~0 (
	.dataa(gnd),
	.datab(out_valid),
	.datac(prev_request_2),
	.datad(top_priority_reg_2),
	.cin(gnd),
	.combout(cout),
	.cout());
defparam \cout~0 .lut_mask = 16'h03FC;
defparam \cout~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sum[1] (
	.dataa(full_addercout_0),
	.datab(top_priority_reg_0),
	.datac(request_1),
	.datad(top_priority_reg_1),
	.cin(gnd),
	.combout(sum_1),
	.cout());
defparam \sum[1] .lut_mask = 16'h2DD2;
defparam \sum[1] .sum_lutc_input = "datac";

cycloneive_lcell_comb \cout~1 (
	.dataa(full_addercout_0),
	.datab(top_priority_reg_2),
	.datac(full_addercout_1),
	.datad(request_2),
	.cin(gnd),
	.combout(cout1),
	.cout());
defparam \cout~1 .lut_mask = 16'h80A8;
defparam \cout~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sum[2] (
	.dataa(out_valid),
	.datab(prev_request_2),
	.datac(top_priority_reg_2),
	.datad(full_addercout_1),
	.cin(gnd),
	.combout(sum_2),
	.cout());
defparam \sum[2] .lut_mask = 16'hE11E;
defparam \sum[2] .sum_lutc_input = "datac";

endmodule

module flashLoader_flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller (
	hold_waitrequest1,
	mem_waitrequest,
	mem_rddata_0,
	mem_rddata_1,
	mem_rddata_2,
	mem_rddata_3,
	mem_rddata_4,
	mem_rddata_5,
	mem_rddata_6,
	mem_rddata_7,
	mem_rddata_8,
	mem_rddata_9,
	mem_rddata_10,
	mem_rddata_11,
	mem_rddata_12,
	mem_rddata_13,
	mem_rddata_14,
	mem_rddata_15,
	mem_rddata_16,
	mem_rddata_17,
	mem_rddata_18,
	mem_rddata_19,
	mem_rddata_20,
	mem_rddata_21,
	mem_rddata_22,
	mem_rddata_23,
	mem_rddata_24,
	mem_rddata_25,
	mem_rddata_26,
	mem_rddata_27,
	mem_rddata_28,
	mem_rddata_29,
	mem_rddata_30,
	mem_rddata_31,
	mem_rddatavalid1,
	csr_wr_inst_data_0,
	csr_rd_inst_data_0,
	altera_reset_synchronizer_int_chain_out,
	csr_wr_inst_data_1,
	csr_rd_inst_data_1,
	csr_wr_inst_data_2,
	csr_rd_inst_data_2,
	csr_wr_inst_data_3,
	csr_rd_inst_data_3,
	csr_wr_inst_data_4,
	csr_rd_inst_data_4,
	csr_wr_inst_data_5,
	csr_rd_inst_data_5,
	csr_wr_inst_data_6,
	csr_rd_inst_data_6,
	csr_wr_inst_data_7,
	csr_rd_inst_data_7,
	csr_rd_inst_data_8,
	csr_control_data_8,
	csr_wr_inst_data_8,
	csr_rd_inst_data_9,
	csr_wr_inst_data_9,
	csr_rd_inst_data_10,
	csr_wr_inst_data_10,
	csr_rd_inst_data_11,
	csr_wr_inst_data_11,
	csr_rd_inst_data_12,
	csr_wr_inst_data_12,
	csr_wr_inst_data_13,
	csr_wr_inst_data_14,
	csr_wr_inst_data_15,
	stateST_SEND_DUMMY_RSP,
	out_valid,
	out_endofpacket,
	out_data_0,
	out_rsp_data_0,
	current_stateSTATE_READ_DATA,
	out_rsp_data_1,
	out_rsp_data_2,
	out_rsp_data_3,
	out_rsp_data_4,
	out_rsp_data_5,
	out_rsp_data_6,
	out_rsp_data_7,
	out_rsp_data_8,
	out_rsp_data_9,
	out_rsp_data_10,
	out_rsp_data_11,
	out_rsp_data_12,
	out_rsp_data_13,
	out_rsp_data_14,
	out_rsp_data_15,
	out_rsp_data_16,
	out_rsp_data_17,
	out_rsp_data_18,
	out_rsp_data_19,
	out_rsp_data_20,
	out_rsp_data_21,
	out_rsp_data_22,
	out_rsp_data_23,
	out_rsp_data_24,
	out_rsp_data_25,
	out_rsp_data_26,
	out_rsp_data_27,
	out_rsp_data_28,
	out_rsp_data_29,
	out_rsp_data_30,
	out_rsp_data_31,
	in_cmd_channel_reg_0,
	saved_grant_0,
	current_stateSTATE_WR_CMD,
	current_stateSTATE_STATUS_CMD,
	current_stateSTATE_POLL_CMD,
	current_stateSTATE_READ_CMD,
	WideOr13,
	current_stateSTATE_WR_DATA,
	cmd_valid,
	Selector18,
	adap_out_cmd_ready,
	Selector181,
	sink0_ready,
	is_burst_reg1,
	mem_write_data_reg_30,
	mem_byteenable_reg_0,
	mem_byteenable_reg_3,
	mem_byteenable_reg_2,
	mem_byteenable_reg_1,
	out_payload_30,
	cmd_valid1,
	mem_write_data_reg_29,
	out_payload_29,
	mem_write_data_reg_28,
	out_payload_28,
	mem_write_data_reg_27,
	out_payload_27,
	out_payload_32,
	cmd_data_11,
	Add1,
	Selector20,
	out_payload_18,
	mem_write_data_reg_18,
	Add11,
	mem_write_data_reg_19,
	out_payload_19,
	mem_write_data_reg_21,
	out_payload_21,
	mem_burstcount_reg_1,
	mem_write_data_reg_20,
	out_payload_20,
	mem_burstcount_reg_0,
	mem_write_data_reg_22,
	out_payload_22,
	mem_burstcount_reg_2,
	mem_write_data_reg_23,
	out_payload_23,
	mem_burstcount_reg_3,
	mem_write_data_reg_24,
	out_payload_24,
	mem_burstcount_reg_4,
	mem_write_data_reg_25,
	out_payload_25,
	mem_burstcount_reg_5,
	mem_write_data_reg_26,
	out_payload_26,
	mem_burstcount_reg_6,
	cmd_data_10,
	cmd_data_8,
	cmd_data_13,
	mem_write_data_reg_17,
	out_payload_17,
	mem_write_data_reg_16,
	out_payload_16,
	mem_write_data_reg_31,
	cmd_data_15,
	cmd_data_14,
	cmd_data_9,
	mem_addr_reg_6,
	mem_addr_reg_14,
	addr_bytes_xip_0,
	out_payload_0,
	cmd_data_0,
	mem_addr_reg_10,
	mem_addr_reg_18,
	mem_addr_reg_2,
	out_payload_4,
	cmd_data_4,
	mem_addr_reg_8,
	mem_addr_reg_16,
	mem_addr_reg_0,
	out_payload_2,
	cmd_data_2,
	mem_addr_reg_15,
	mem_addr_reg_7,
	WideOr19,
	out_payload_1,
	cmd_data_1,
	mem_addr_reg_17,
	mem_addr_reg_9,
	mem_addr_reg_1,
	out_payload_3,
	cmd_data_3,
	mem_addr_reg_19,
	mem_addr_reg_11,
	mem_addr_reg_3,
	out_payload_5,
	cmd_data_5,
	mem_addr_reg_12,
	mem_addr_reg_20,
	mem_addr_reg_4,
	out_payload_6,
	cmd_data_6,
	mem_addr_reg_13,
	mem_addr_reg_5,
	out_payload_7,
	cmd_data_7,
	cmd_data_12,
	out_payload_31,
	clk_clk,
	avl_mem_read,
	mem_burstcount,
	avl_mem_write,
	avl_mem_byteenable_0,
	avl_mem_byteenable_1,
	avl_mem_byteenable_2,
	avl_mem_byteenable_3,
	avl_mem_writedata_30,
	avl_mem_writedata_29,
	avl_mem_writedata_28,
	avl_mem_writedata_27,
	avl_mem_writedata_11,
	avl_mem_writedata_18,
	avl_mem_writedata_19,
	avl_mem_writedata_21,
	avl_mem_writedata_20,
	avl_mem_writedata_22,
	avl_mem_writedata_23,
	avl_mem_writedata_24,
	avl_mem_writedata_25,
	avl_mem_writedata_26,
	avl_mem_writedata_10,
	avl_mem_writedata_8,
	avl_mem_writedata_13,
	avl_mem_writedata_17,
	avl_mem_writedata_16,
	avl_mem_writedata_15,
	avl_mem_writedata_31,
	avl_mem_writedata_14,
	avl_mem_writedata_9,
	mem_addr,
	avl_mem_writedata_0,
	avl_mem_writedata_4,
	avl_mem_writedata_12,
	avl_mem_writedata_2,
	avl_mem_writedata_1,
	avl_mem_writedata_3,
	avl_mem_writedata_5,
	avl_mem_writedata_6,
	avl_mem_writedata_7)/* synthesis synthesis_greybox=0 */;
output 	hold_waitrequest1;
output 	mem_waitrequest;
output 	mem_rddata_0;
output 	mem_rddata_1;
output 	mem_rddata_2;
output 	mem_rddata_3;
output 	mem_rddata_4;
output 	mem_rddata_5;
output 	mem_rddata_6;
output 	mem_rddata_7;
output 	mem_rddata_8;
output 	mem_rddata_9;
output 	mem_rddata_10;
output 	mem_rddata_11;
output 	mem_rddata_12;
output 	mem_rddata_13;
output 	mem_rddata_14;
output 	mem_rddata_15;
output 	mem_rddata_16;
output 	mem_rddata_17;
output 	mem_rddata_18;
output 	mem_rddata_19;
output 	mem_rddata_20;
output 	mem_rddata_21;
output 	mem_rddata_22;
output 	mem_rddata_23;
output 	mem_rddata_24;
output 	mem_rddata_25;
output 	mem_rddata_26;
output 	mem_rddata_27;
output 	mem_rddata_28;
output 	mem_rddata_29;
output 	mem_rddata_30;
output 	mem_rddata_31;
output 	mem_rddatavalid1;
input 	csr_wr_inst_data_0;
input 	csr_rd_inst_data_0;
input 	altera_reset_synchronizer_int_chain_out;
input 	csr_wr_inst_data_1;
input 	csr_rd_inst_data_1;
input 	csr_wr_inst_data_2;
input 	csr_rd_inst_data_2;
input 	csr_wr_inst_data_3;
input 	csr_rd_inst_data_3;
input 	csr_wr_inst_data_4;
input 	csr_rd_inst_data_4;
input 	csr_wr_inst_data_5;
input 	csr_rd_inst_data_5;
input 	csr_wr_inst_data_6;
input 	csr_rd_inst_data_6;
input 	csr_wr_inst_data_7;
input 	csr_rd_inst_data_7;
input 	csr_rd_inst_data_8;
input 	csr_control_data_8;
input 	csr_wr_inst_data_8;
input 	csr_rd_inst_data_9;
input 	csr_wr_inst_data_9;
input 	csr_rd_inst_data_10;
input 	csr_wr_inst_data_10;
input 	csr_rd_inst_data_11;
input 	csr_wr_inst_data_11;
input 	csr_rd_inst_data_12;
input 	csr_wr_inst_data_12;
input 	csr_wr_inst_data_13;
input 	csr_wr_inst_data_14;
input 	csr_wr_inst_data_15;
input 	stateST_SEND_DUMMY_RSP;
input 	out_valid;
input 	out_endofpacket;
input 	out_data_0;
input 	out_rsp_data_0;
output 	current_stateSTATE_READ_DATA;
input 	out_rsp_data_1;
input 	out_rsp_data_2;
input 	out_rsp_data_3;
input 	out_rsp_data_4;
input 	out_rsp_data_5;
input 	out_rsp_data_6;
input 	out_rsp_data_7;
input 	out_rsp_data_8;
input 	out_rsp_data_9;
input 	out_rsp_data_10;
input 	out_rsp_data_11;
input 	out_rsp_data_12;
input 	out_rsp_data_13;
input 	out_rsp_data_14;
input 	out_rsp_data_15;
input 	out_rsp_data_16;
input 	out_rsp_data_17;
input 	out_rsp_data_18;
input 	out_rsp_data_19;
input 	out_rsp_data_20;
input 	out_rsp_data_21;
input 	out_rsp_data_22;
input 	out_rsp_data_23;
input 	out_rsp_data_24;
input 	out_rsp_data_25;
input 	out_rsp_data_26;
input 	out_rsp_data_27;
input 	out_rsp_data_28;
input 	out_rsp_data_29;
input 	out_rsp_data_30;
input 	out_rsp_data_31;
input 	in_cmd_channel_reg_0;
input 	saved_grant_0;
output 	current_stateSTATE_WR_CMD;
output 	current_stateSTATE_STATUS_CMD;
output 	current_stateSTATE_POLL_CMD;
output 	current_stateSTATE_READ_CMD;
output 	WideOr13;
output 	current_stateSTATE_WR_DATA;
output 	cmd_valid;
input 	Selector18;
input 	adap_out_cmd_ready;
input 	Selector181;
input 	sink0_ready;
output 	is_burst_reg1;
output 	mem_write_data_reg_30;
output 	mem_byteenable_reg_0;
output 	mem_byteenable_reg_3;
output 	mem_byteenable_reg_2;
output 	mem_byteenable_reg_1;
output 	out_payload_30;
output 	cmd_valid1;
output 	mem_write_data_reg_29;
output 	out_payload_29;
output 	mem_write_data_reg_28;
output 	out_payload_28;
output 	mem_write_data_reg_27;
output 	out_payload_27;
output 	out_payload_32;
output 	cmd_data_11;
output 	Add1;
output 	Selector20;
output 	out_payload_18;
output 	mem_write_data_reg_18;
output 	Add11;
output 	mem_write_data_reg_19;
output 	out_payload_19;
output 	mem_write_data_reg_21;
output 	out_payload_21;
output 	mem_burstcount_reg_1;
output 	mem_write_data_reg_20;
output 	out_payload_20;
output 	mem_burstcount_reg_0;
output 	mem_write_data_reg_22;
output 	out_payload_22;
output 	mem_burstcount_reg_2;
output 	mem_write_data_reg_23;
output 	out_payload_23;
output 	mem_burstcount_reg_3;
output 	mem_write_data_reg_24;
output 	out_payload_24;
output 	mem_burstcount_reg_4;
output 	mem_write_data_reg_25;
output 	out_payload_25;
output 	mem_burstcount_reg_5;
output 	mem_write_data_reg_26;
output 	out_payload_26;
output 	mem_burstcount_reg_6;
output 	cmd_data_10;
output 	cmd_data_8;
output 	cmd_data_13;
output 	mem_write_data_reg_17;
output 	out_payload_17;
output 	mem_write_data_reg_16;
output 	out_payload_16;
output 	mem_write_data_reg_31;
output 	cmd_data_15;
output 	cmd_data_14;
output 	cmd_data_9;
output 	mem_addr_reg_6;
output 	mem_addr_reg_14;
output 	addr_bytes_xip_0;
output 	out_payload_0;
output 	cmd_data_0;
output 	mem_addr_reg_10;
output 	mem_addr_reg_18;
output 	mem_addr_reg_2;
output 	out_payload_4;
output 	cmd_data_4;
output 	mem_addr_reg_8;
output 	mem_addr_reg_16;
output 	mem_addr_reg_0;
output 	out_payload_2;
output 	cmd_data_2;
output 	mem_addr_reg_15;
output 	mem_addr_reg_7;
output 	WideOr19;
output 	out_payload_1;
output 	cmd_data_1;
output 	mem_addr_reg_17;
output 	mem_addr_reg_9;
output 	mem_addr_reg_1;
output 	out_payload_3;
output 	cmd_data_3;
output 	mem_addr_reg_19;
output 	mem_addr_reg_11;
output 	mem_addr_reg_3;
output 	out_payload_5;
output 	cmd_data_5;
output 	mem_addr_reg_12;
output 	mem_addr_reg_20;
output 	mem_addr_reg_4;
output 	out_payload_6;
output 	cmd_data_6;
output 	mem_addr_reg_13;
output 	mem_addr_reg_5;
output 	out_payload_7;
output 	cmd_data_7;
output 	cmd_data_12;
output 	out_payload_31;
input 	clk_clk;
input 	avl_mem_read;
input 	[6:0] mem_burstcount;
input 	avl_mem_write;
input 	avl_mem_byteenable_0;
input 	avl_mem_byteenable_1;
input 	avl_mem_byteenable_2;
input 	avl_mem_byteenable_3;
input 	avl_mem_writedata_30;
input 	avl_mem_writedata_29;
input 	avl_mem_writedata_28;
input 	avl_mem_writedata_27;
input 	avl_mem_writedata_11;
input 	avl_mem_writedata_18;
input 	avl_mem_writedata_19;
input 	avl_mem_writedata_21;
input 	avl_mem_writedata_20;
input 	avl_mem_writedata_22;
input 	avl_mem_writedata_23;
input 	avl_mem_writedata_24;
input 	avl_mem_writedata_25;
input 	avl_mem_writedata_26;
input 	avl_mem_writedata_10;
input 	avl_mem_writedata_8;
input 	avl_mem_writedata_13;
input 	avl_mem_writedata_17;
input 	avl_mem_writedata_16;
input 	avl_mem_writedata_15;
input 	avl_mem_writedata_31;
input 	avl_mem_writedata_14;
input 	avl_mem_writedata_9;
input 	[31:0] mem_addr;
input 	avl_mem_writedata_0;
input 	avl_mem_writedata_4;
input 	avl_mem_writedata_12;
input 	avl_mem_writedata_2;
input 	avl_mem_writedata_1;
input 	avl_mem_writedata_3;
input 	avl_mem_writedata_5;
input 	avl_mem_writedata_6;
input 	avl_mem_writedata_7;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \avst_fifo_inst|avst_fifo|full~q ;
wire \avst_fifo_inst|avst_fifo|out_valid~q ;
wire \avst_fifo_inst|avst_fifo|out_payload[11]~q ;
wire \avst_fifo_inst|avst_fifo|out_payload[10]~q ;
wire \avst_fifo_inst|avst_fifo|out_payload[8]~q ;
wire \avst_fifo_inst|avst_fifo|out_payload[13]~q ;
wire \avst_fifo_inst|avst_fifo|out_payload[15]~q ;
wire \avst_fifo_inst|avst_fifo|out_payload[14]~q ;
wire \avst_fifo_inst|avst_fifo|out_payload[9]~q ;
wire \avst_fifo_inst|avst_fifo|out_payload[12]~q ;
wire \always0~0_combout ;
wire \Selector8~0_combout ;
wire \current_state.STATE_POLL_RSP~q ;
wire \Equal3~0_combout ;
wire \Equal3~1_combout ;
wire \busy~0_combout ;
wire \Selector12~0_combout ;
wire \current_state.STATE_COMPLETE~q ;
wire \burstcount_register[0]~7_combout ;
wire \Equal0~0_combout ;
wire \sop_enable~0_combout ;
wire \mem_wr_combi~0_combout ;
wire \sop_enable~q ;
wire \burstcount_register~9_combout ;
wire \burstcount_register[0]~q ;
wire \internal_burstcount[0]~0_combout ;
wire \burstcount_register[0]~8 ;
wire \burstcount_register[1]~10_combout ;
wire \burstcount_register[1]~q ;
wire \internal_burstcount[1]~3_combout ;
wire \burstcount_register[1]~11 ;
wire \burstcount_register[2]~12_combout ;
wire \burstcount_register[2]~q ;
wire \internal_burstcount[2]~2_combout ;
wire \burstcount_register[2]~13 ;
wire \burstcount_register[3]~14_combout ;
wire \burstcount_register[3]~q ;
wire \internal_burstcount[3]~6_combout ;
wire \burstcount_register[3]~15 ;
wire \burstcount_register[4]~16_combout ;
wire \burstcount_register[4]~q ;
wire \internal_burstcount[4]~5_combout ;
wire \burstcount_register[4]~17 ;
wire \burstcount_register[5]~18_combout ;
wire \burstcount_register[5]~q ;
wire \internal_burstcount[5]~4_combout ;
wire \burstcount_register[5]~19 ;
wire \burstcount_register[6]~20_combout ;
wire \burstcount_register[6]~q ;
wire \internal_burstcount[6]~1_combout ;
wire \Equal2~0_combout ;
wire \Equal2~1_combout ;
wire \Selector0~0_combout ;
wire \Selector0~1_combout ;
wire \Selector0~2_combout ;
wire \current_state.STATE_IDLE~q ;
wire \mem_rddatavalid~0_combout ;
wire \Selector11~0_combout ;
wire \Selector2~0_combout ;
wire \current_state.STATE_STATUS_RSP~q ;
wire \Selector3~0_combout ;
wire \Selector3~1_combout ;
wire \current_state.STATE_WRENABLE_CMD~q ;
wire \Selector4~0_combout ;
wire \current_state.STATE_WRENABLE_RSP~q ;
wire \Selector5~0_combout ;
wire \next_state~0_combout ;
wire \Selector1~0_combout ;
wire \fifo_in_valid~0_combout ;
wire \Selector10~0_combout ;
wire \Selector1~1_combout ;
wire \Selector1~2_combout ;
wire \Selector7~0_combout ;
wire \Selector7~1_combout ;
wire \Selector10~1_combout ;
wire \Selector6~0_combout ;
wire \always10~2_combout ;
wire \mem_byteenable_reg[0]~0_combout ;
wire \mem_byteenable_reg[0]~1_combout ;
wire \is_burst_reg~0_combout ;
wire \mem_byteenable_reg~2_combout ;
wire \mem_byteenable_reg[0]~3_combout ;
wire \mem_byteenable_reg~4_combout ;
wire \mem_byteenable_reg~5_combout ;
wire \mem_byteenable_reg~6_combout ;
wire \mem_write_data_reg[11]~q ;
wire \cmd_data[11]~4_combout ;
wire \Add1~0_combout ;
wire \cmd_data[8]~5_combout ;
wire \cmd_data[8]~88_combout ;
wire \Selector17~0_combout ;
wire \cmd_data[8]~6_combout ;
wire \cmd_data[11]~7_combout ;
wire \mem_write_data_reg[10]~q ;
wire \cmd_data[10]~8_combout ;
wire \cmd_data[10]~9_combout ;
wire \mem_write_data_reg[8]~q ;
wire \cmd_data[8]~10_combout ;
wire \cmd_data[8]~11_combout ;
wire \mem_write_data_reg[13]~q ;
wire \cmd_data[13]~12_combout ;
wire \Selector15~0_combout ;
wire \cmd_data[13]~13_combout ;
wire \mem_write_data_reg[15]~q ;
wire \cmd_data[15]~14_combout ;
wire \cmd_data[14]~15_combout ;
wire \cmd_data[14]~89_combout ;
wire \cmd_data[15]~16_combout ;
wire \cmd_data[15]~17_combout ;
wire \mem_write_data_reg[14]~q ;
wire \cmd_data[14]~18_combout ;
wire \cmd_data[14]~19_combout ;
wire \cmd_data[14]~20_combout ;
wire \mem_write_data_reg[9]~q ;
wire \cmd_data[9]~21_combout ;
wire \Selector19~0_combout ;
wire \cmd_data[9]~22_combout ;
wire \cmd_data[0]~23_combout ;
wire \cmd_data[2]~24_combout ;
wire \cmd_data[2]~25_combout ;
wire \mem_write_data_reg[0]~q ;
wire \cmd_data[2]~26_combout ;
wire \cmd_data[0]~27_combout ;
wire \cmd_data[2]~28_combout ;
wire \cmd_data[0]~29_combout ;
wire \cmd_data[0]~30_combout ;
wire \cmd_data[0]~31_combout ;
wire \cmd_data[2]~32_combout ;
wire \cmd_data[2]~33_combout ;
wire \cmd_data[2]~34_combout ;
wire \cmd_data[0]~35_combout ;
wire \cmd_data[4]~37_combout ;
wire \mem_write_data_reg[4]~q ;
wire \cmd_data[4]~38_combout ;
wire \mem_write_data_reg[12]~q ;
wire \cmd_data[4]~39_combout ;
wire \cmd_data[4]~40_combout ;
wire \cmd_data[4]~41_combout ;
wire \cmd_data[4]~42_combout ;
wire \cmd_data[2]~44_combout ;
wire \mem_write_data_reg[2]~q ;
wire \cmd_data[2]~45_combout ;
wire \cmd_data[2]~46_combout ;
wire \cmd_data[2]~47_combout ;
wire \cmd_data[2]~48_combout ;
wire \cmd_data[2]~49_combout ;
wire \cmd_data[1]~51_combout ;
wire \mem_write_data_reg[1]~q ;
wire \cmd_data[1]~52_combout ;
wire \cmd_data[1]~53_combout ;
wire \cmd_data[1]~54_combout ;
wire \cmd_data[1]~55_combout ;
wire \cmd_data[1]~56_combout ;
wire \cmd_data[3]~58_combout ;
wire \mem_write_data_reg[3]~q ;
wire \cmd_data[3]~59_combout ;
wire \cmd_data[3]~60_combout ;
wire \cmd_data[3]~61_combout ;
wire \cmd_data[3]~62_combout ;
wire \cmd_data[3]~63_combout ;
wire \cmd_data[5]~65_combout ;
wire \mem_write_data_reg[5]~q ;
wire \cmd_data[5]~66_combout ;
wire \cmd_data[5]~67_combout ;
wire \cmd_data[5]~68_combout ;
wire \cmd_data[5]~69_combout ;
wire \cmd_data[5]~70_combout ;
wire \cmd_data[6]~72_combout ;
wire \mem_write_data_reg[6]~q ;
wire \cmd_data[6]~73_combout ;
wire \cmd_data[6]~74_combout ;
wire \cmd_data[6]~75_combout ;
wire \cmd_data[6]~76_combout ;
wire \cmd_data[6]~77_combout ;
wire \cmd_data[7]~79_combout ;
wire \mem_write_data_reg[7]~q ;
wire \cmd_data[7]~80_combout ;
wire \cmd_data[7]~81_combout ;
wire \cmd_data[7]~82_combout ;
wire \cmd_data[7]~83_combout ;
wire \cmd_data[7]~84_combout ;
wire \cmd_data[12]~86_combout ;
wire \Selector16~0_combout ;
wire \Selector16~1_combout ;
wire \cmd_data[12]~87_combout ;


flashLoader_avst_fifo avst_fifo_inst(
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.Equal2(\Equal2~1_combout ),
	.full(\avst_fifo_inst|avst_fifo|full~q ),
	.saved_grant_0(saved_grant_0),
	.out_valid(\avst_fifo_inst|avst_fifo|out_valid~q ),
	.current_stateSTATE_WR_DATA(current_stateSTATE_WR_DATA),
	.Selector18(Selector18),
	.adap_out_cmd_ready(adap_out_cmd_ready),
	.Selector181(Selector181),
	.mem_wr_combi(\mem_wr_combi~0_combout ),
	.sink0_ready(sink0_ready),
	.out_payload_30(out_payload_30),
	.out_payload_29(out_payload_29),
	.out_payload_28(out_payload_28),
	.out_payload_27(out_payload_27),
	.out_payload_32(out_payload_32),
	.fifo_in_valid(\fifo_in_valid~0_combout ),
	.out_payload_11(\avst_fifo_inst|avst_fifo|out_payload[11]~q ),
	.out_payload_18(out_payload_18),
	.out_payload_19(out_payload_19),
	.out_payload_21(out_payload_21),
	.out_payload_20(out_payload_20),
	.out_payload_22(out_payload_22),
	.out_payload_23(out_payload_23),
	.out_payload_24(out_payload_24),
	.out_payload_25(out_payload_25),
	.out_payload_26(out_payload_26),
	.out_payload_10(\avst_fifo_inst|avst_fifo|out_payload[10]~q ),
	.out_payload_8(\avst_fifo_inst|avst_fifo|out_payload[8]~q ),
	.out_payload_13(\avst_fifo_inst|avst_fifo|out_payload[13]~q ),
	.out_payload_17(out_payload_17),
	.out_payload_16(out_payload_16),
	.out_payload_15(\avst_fifo_inst|avst_fifo|out_payload[15]~q ),
	.out_payload_14(\avst_fifo_inst|avst_fifo|out_payload[14]~q ),
	.out_payload_9(\avst_fifo_inst|avst_fifo|out_payload[9]~q ),
	.out_payload_0(out_payload_0),
	.out_payload_4(out_payload_4),
	.out_payload_2(out_payload_2),
	.out_payload_1(out_payload_1),
	.out_payload_3(out_payload_3),
	.out_payload_5(out_payload_5),
	.out_payload_6(out_payload_6),
	.out_payload_7(out_payload_7),
	.out_payload_12(\avst_fifo_inst|avst_fifo|out_payload[12]~q ),
	.out_payload_31(out_payload_31),
	.clk_clk(clk_clk),
	.avl_mem_writedata_30(avl_mem_writedata_30),
	.avl_mem_writedata_29(avl_mem_writedata_29),
	.avl_mem_writedata_28(avl_mem_writedata_28),
	.avl_mem_writedata_27(avl_mem_writedata_27),
	.avl_mem_writedata_11(avl_mem_writedata_11),
	.avl_mem_writedata_18(avl_mem_writedata_18),
	.avl_mem_writedata_19(avl_mem_writedata_19),
	.avl_mem_writedata_21(avl_mem_writedata_21),
	.avl_mem_writedata_20(avl_mem_writedata_20),
	.avl_mem_writedata_22(avl_mem_writedata_22),
	.avl_mem_writedata_23(avl_mem_writedata_23),
	.avl_mem_writedata_24(avl_mem_writedata_24),
	.avl_mem_writedata_25(avl_mem_writedata_25),
	.avl_mem_writedata_26(avl_mem_writedata_26),
	.avl_mem_writedata_10(avl_mem_writedata_10),
	.avl_mem_writedata_8(avl_mem_writedata_8),
	.avl_mem_writedata_13(avl_mem_writedata_13),
	.avl_mem_writedata_17(avl_mem_writedata_17),
	.avl_mem_writedata_16(avl_mem_writedata_16),
	.avl_mem_writedata_15(avl_mem_writedata_15),
	.avl_mem_writedata_31(avl_mem_writedata_31),
	.avl_mem_writedata_14(avl_mem_writedata_14),
	.avl_mem_writedata_9(avl_mem_writedata_9),
	.avl_mem_writedata_0(avl_mem_writedata_0),
	.avl_mem_writedata_4(avl_mem_writedata_4),
	.avl_mem_writedata_12(avl_mem_writedata_12),
	.avl_mem_writedata_2(avl_mem_writedata_2),
	.avl_mem_writedata_1(avl_mem_writedata_1),
	.avl_mem_writedata_3(avl_mem_writedata_3),
	.avl_mem_writedata_5(avl_mem_writedata_5),
	.avl_mem_writedata_6(avl_mem_writedata_6),
	.avl_mem_writedata_7(avl_mem_writedata_7));

dffeas hold_waitrequest(
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(hold_waitrequest1),
	.prn(vcc));
defparam hold_waitrequest.is_wysiwyg = "true";
defparam hold_waitrequest.power_up = "low";

cycloneive_lcell_comb \mem_waitrequest~0 (
	.dataa(hold_waitrequest1),
	.datab(gnd),
	.datac(gnd),
	.datad(\current_state.STATE_IDLE~q ),
	.cin(gnd),
	.combout(mem_waitrequest),
	.cout());
defparam \mem_waitrequest~0 .lut_mask = 16'h00AA;
defparam \mem_waitrequest~0 .sum_lutc_input = "datac";

dffeas \mem_rddata[0] (
	.clk(clk_clk),
	.d(out_rsp_data_0),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_0),
	.prn(vcc));
defparam \mem_rddata[0] .is_wysiwyg = "true";
defparam \mem_rddata[0] .power_up = "low";

dffeas \mem_rddata[1] (
	.clk(clk_clk),
	.d(out_rsp_data_1),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_1),
	.prn(vcc));
defparam \mem_rddata[1] .is_wysiwyg = "true";
defparam \mem_rddata[1] .power_up = "low";

dffeas \mem_rddata[2] (
	.clk(clk_clk),
	.d(out_rsp_data_2),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_2),
	.prn(vcc));
defparam \mem_rddata[2] .is_wysiwyg = "true";
defparam \mem_rddata[2] .power_up = "low";

dffeas \mem_rddata[3] (
	.clk(clk_clk),
	.d(out_rsp_data_3),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_3),
	.prn(vcc));
defparam \mem_rddata[3] .is_wysiwyg = "true";
defparam \mem_rddata[3] .power_up = "low";

dffeas \mem_rddata[4] (
	.clk(clk_clk),
	.d(out_rsp_data_4),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_4),
	.prn(vcc));
defparam \mem_rddata[4] .is_wysiwyg = "true";
defparam \mem_rddata[4] .power_up = "low";

dffeas \mem_rddata[5] (
	.clk(clk_clk),
	.d(out_rsp_data_5),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_5),
	.prn(vcc));
defparam \mem_rddata[5] .is_wysiwyg = "true";
defparam \mem_rddata[5] .power_up = "low";

dffeas \mem_rddata[6] (
	.clk(clk_clk),
	.d(out_rsp_data_6),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_6),
	.prn(vcc));
defparam \mem_rddata[6] .is_wysiwyg = "true";
defparam \mem_rddata[6] .power_up = "low";

dffeas \mem_rddata[7] (
	.clk(clk_clk),
	.d(out_rsp_data_7),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_7),
	.prn(vcc));
defparam \mem_rddata[7] .is_wysiwyg = "true";
defparam \mem_rddata[7] .power_up = "low";

dffeas \mem_rddata[8] (
	.clk(clk_clk),
	.d(out_rsp_data_8),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_8),
	.prn(vcc));
defparam \mem_rddata[8] .is_wysiwyg = "true";
defparam \mem_rddata[8] .power_up = "low";

dffeas \mem_rddata[9] (
	.clk(clk_clk),
	.d(out_rsp_data_9),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_9),
	.prn(vcc));
defparam \mem_rddata[9] .is_wysiwyg = "true";
defparam \mem_rddata[9] .power_up = "low";

dffeas \mem_rddata[10] (
	.clk(clk_clk),
	.d(out_rsp_data_10),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_10),
	.prn(vcc));
defparam \mem_rddata[10] .is_wysiwyg = "true";
defparam \mem_rddata[10] .power_up = "low";

dffeas \mem_rddata[11] (
	.clk(clk_clk),
	.d(out_rsp_data_11),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_11),
	.prn(vcc));
defparam \mem_rddata[11] .is_wysiwyg = "true";
defparam \mem_rddata[11] .power_up = "low";

dffeas \mem_rddata[12] (
	.clk(clk_clk),
	.d(out_rsp_data_12),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_12),
	.prn(vcc));
defparam \mem_rddata[12] .is_wysiwyg = "true";
defparam \mem_rddata[12] .power_up = "low";

dffeas \mem_rddata[13] (
	.clk(clk_clk),
	.d(out_rsp_data_13),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_13),
	.prn(vcc));
defparam \mem_rddata[13] .is_wysiwyg = "true";
defparam \mem_rddata[13] .power_up = "low";

dffeas \mem_rddata[14] (
	.clk(clk_clk),
	.d(out_rsp_data_14),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_14),
	.prn(vcc));
defparam \mem_rddata[14] .is_wysiwyg = "true";
defparam \mem_rddata[14] .power_up = "low";

dffeas \mem_rddata[15] (
	.clk(clk_clk),
	.d(out_rsp_data_15),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_15),
	.prn(vcc));
defparam \mem_rddata[15] .is_wysiwyg = "true";
defparam \mem_rddata[15] .power_up = "low";

dffeas \mem_rddata[16] (
	.clk(clk_clk),
	.d(out_rsp_data_16),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_16),
	.prn(vcc));
defparam \mem_rddata[16] .is_wysiwyg = "true";
defparam \mem_rddata[16] .power_up = "low";

dffeas \mem_rddata[17] (
	.clk(clk_clk),
	.d(out_rsp_data_17),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_17),
	.prn(vcc));
defparam \mem_rddata[17] .is_wysiwyg = "true";
defparam \mem_rddata[17] .power_up = "low";

dffeas \mem_rddata[18] (
	.clk(clk_clk),
	.d(out_rsp_data_18),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_18),
	.prn(vcc));
defparam \mem_rddata[18] .is_wysiwyg = "true";
defparam \mem_rddata[18] .power_up = "low";

dffeas \mem_rddata[19] (
	.clk(clk_clk),
	.d(out_rsp_data_19),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_19),
	.prn(vcc));
defparam \mem_rddata[19] .is_wysiwyg = "true";
defparam \mem_rddata[19] .power_up = "low";

dffeas \mem_rddata[20] (
	.clk(clk_clk),
	.d(out_rsp_data_20),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_20),
	.prn(vcc));
defparam \mem_rddata[20] .is_wysiwyg = "true";
defparam \mem_rddata[20] .power_up = "low";

dffeas \mem_rddata[21] (
	.clk(clk_clk),
	.d(out_rsp_data_21),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_21),
	.prn(vcc));
defparam \mem_rddata[21] .is_wysiwyg = "true";
defparam \mem_rddata[21] .power_up = "low";

dffeas \mem_rddata[22] (
	.clk(clk_clk),
	.d(out_rsp_data_22),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_22),
	.prn(vcc));
defparam \mem_rddata[22] .is_wysiwyg = "true";
defparam \mem_rddata[22] .power_up = "low";

dffeas \mem_rddata[23] (
	.clk(clk_clk),
	.d(out_rsp_data_23),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_23),
	.prn(vcc));
defparam \mem_rddata[23] .is_wysiwyg = "true";
defparam \mem_rddata[23] .power_up = "low";

dffeas \mem_rddata[24] (
	.clk(clk_clk),
	.d(out_rsp_data_24),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_24),
	.prn(vcc));
defparam \mem_rddata[24] .is_wysiwyg = "true";
defparam \mem_rddata[24] .power_up = "low";

dffeas \mem_rddata[25] (
	.clk(clk_clk),
	.d(out_rsp_data_25),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_25),
	.prn(vcc));
defparam \mem_rddata[25] .is_wysiwyg = "true";
defparam \mem_rddata[25] .power_up = "low";

dffeas \mem_rddata[26] (
	.clk(clk_clk),
	.d(out_rsp_data_26),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_26),
	.prn(vcc));
defparam \mem_rddata[26] .is_wysiwyg = "true";
defparam \mem_rddata[26] .power_up = "low";

dffeas \mem_rddata[27] (
	.clk(clk_clk),
	.d(out_rsp_data_27),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_27),
	.prn(vcc));
defparam \mem_rddata[27] .is_wysiwyg = "true";
defparam \mem_rddata[27] .power_up = "low";

dffeas \mem_rddata[28] (
	.clk(clk_clk),
	.d(out_rsp_data_28),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_28),
	.prn(vcc));
defparam \mem_rddata[28] .is_wysiwyg = "true";
defparam \mem_rddata[28] .power_up = "low";

dffeas \mem_rddata[29] (
	.clk(clk_clk),
	.d(out_rsp_data_29),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_29),
	.prn(vcc));
defparam \mem_rddata[29] .is_wysiwyg = "true";
defparam \mem_rddata[29] .power_up = "low";

dffeas \mem_rddata[30] (
	.clk(clk_clk),
	.d(out_rsp_data_30),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_30),
	.prn(vcc));
defparam \mem_rddata[30] .is_wysiwyg = "true";
defparam \mem_rddata[30] .power_up = "low";

dffeas \mem_rddata[31] (
	.clk(clk_clk),
	.d(out_rsp_data_31),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(current_stateSTATE_READ_DATA),
	.q(mem_rddata_31),
	.prn(vcc));
defparam \mem_rddata[31] .is_wysiwyg = "true";
defparam \mem_rddata[31] .power_up = "low";

dffeas mem_rddatavalid(
	.clk(clk_clk),
	.d(\mem_rddatavalid~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_rddatavalid1),
	.prn(vcc));
defparam mem_rddatavalid.is_wysiwyg = "true";
defparam mem_rddatavalid.power_up = "low";

dffeas \current_state.STATE_READ_DATA (
	.clk(clk_clk),
	.d(\Selector11~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(current_stateSTATE_READ_DATA),
	.prn(vcc));
defparam \current_state.STATE_READ_DATA .is_wysiwyg = "true";
defparam \current_state.STATE_READ_DATA .power_up = "low";

dffeas \current_state.STATE_WR_CMD (
	.clk(clk_clk),
	.d(\Selector5~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(current_stateSTATE_WR_CMD),
	.prn(vcc));
defparam \current_state.STATE_WR_CMD .is_wysiwyg = "true";
defparam \current_state.STATE_WR_CMD .power_up = "low";

dffeas \current_state.STATE_STATUS_CMD (
	.clk(clk_clk),
	.d(\Selector1~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(current_stateSTATE_STATUS_CMD),
	.prn(vcc));
defparam \current_state.STATE_STATUS_CMD .is_wysiwyg = "true";
defparam \current_state.STATE_STATUS_CMD .power_up = "low";

dffeas \current_state.STATE_POLL_CMD (
	.clk(clk_clk),
	.d(\Selector7~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(current_stateSTATE_POLL_CMD),
	.prn(vcc));
defparam \current_state.STATE_POLL_CMD .is_wysiwyg = "true";
defparam \current_state.STATE_POLL_CMD .power_up = "low";

dffeas \current_state.STATE_READ_CMD (
	.clk(clk_clk),
	.d(\Selector10~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(current_stateSTATE_READ_CMD),
	.prn(vcc));
defparam \current_state.STATE_READ_CMD .is_wysiwyg = "true";
defparam \current_state.STATE_READ_CMD .power_up = "low";

cycloneive_lcell_comb \WideOr13~0 (
	.dataa(current_stateSTATE_STATUS_CMD),
	.datab(\current_state.STATE_WRENABLE_CMD~q ),
	.datac(current_stateSTATE_POLL_CMD),
	.datad(current_stateSTATE_READ_CMD),
	.cin(gnd),
	.combout(WideOr13),
	.cout());
defparam \WideOr13~0 .lut_mask = 16'h0001;
defparam \WideOr13~0 .sum_lutc_input = "datac";

dffeas \current_state.STATE_WR_DATA (
	.clk(clk_clk),
	.d(\Selector6~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(current_stateSTATE_WR_DATA),
	.prn(vcc));
defparam \current_state.STATE_WR_DATA .is_wysiwyg = "true";
defparam \current_state.STATE_WR_DATA .power_up = "low";

cycloneive_lcell_comb \cmd_valid~0 (
	.dataa(\avst_fifo_inst|avst_fifo|out_valid~q ),
	.datab(current_stateSTATE_WR_CMD),
	.datac(WideOr13),
	.datad(current_stateSTATE_WR_DATA),
	.cin(gnd),
	.combout(cmd_valid),
	.cout());
defparam \cmd_valid~0 .lut_mask = 16'hAACF;
defparam \cmd_valid~0 .sum_lutc_input = "datac";

dffeas is_burst_reg(
	.clk(clk_clk),
	.d(\is_burst_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(is_burst_reg1),
	.prn(vcc));
defparam is_burst_reg.is_wysiwyg = "true";
defparam is_burst_reg.power_up = "low";

dffeas \mem_write_data_reg[30] (
	.clk(clk_clk),
	.d(avl_mem_writedata_30),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(mem_write_data_reg_30),
	.prn(vcc));
defparam \mem_write_data_reg[30] .is_wysiwyg = "true";
defparam \mem_write_data_reg[30] .power_up = "low";

dffeas \mem_byteenable_reg[0] (
	.clk(clk_clk),
	.d(\mem_byteenable_reg~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_byteenable_reg_0),
	.prn(vcc));
defparam \mem_byteenable_reg[0] .is_wysiwyg = "true";
defparam \mem_byteenable_reg[0] .power_up = "low";

dffeas \mem_byteenable_reg[3] (
	.clk(clk_clk),
	.d(\mem_byteenable_reg~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_byteenable_reg_3),
	.prn(vcc));
defparam \mem_byteenable_reg[3] .is_wysiwyg = "true";
defparam \mem_byteenable_reg[3] .power_up = "low";

dffeas \mem_byteenable_reg[2] (
	.clk(clk_clk),
	.d(\mem_byteenable_reg~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_byteenable_reg_2),
	.prn(vcc));
defparam \mem_byteenable_reg[2] .is_wysiwyg = "true";
defparam \mem_byteenable_reg[2] .power_up = "low";

dffeas \mem_byteenable_reg[1] (
	.clk(clk_clk),
	.d(\mem_byteenable_reg~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_byteenable_reg_1),
	.prn(vcc));
defparam \mem_byteenable_reg[1] .is_wysiwyg = "true";
defparam \mem_byteenable_reg[1] .power_up = "low";

cycloneive_lcell_comb \cmd_valid~1 (
	.dataa(current_stateSTATE_WR_CMD),
	.datab(gnd),
	.datac(WideOr13),
	.datad(current_stateSTATE_WR_DATA),
	.cin(gnd),
	.combout(cmd_valid1),
	.cout());
defparam \cmd_valid~1 .lut_mask = 16'h00AF;
defparam \cmd_valid~1 .sum_lutc_input = "datac";

dffeas \mem_write_data_reg[29] (
	.clk(clk_clk),
	.d(avl_mem_writedata_29),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(mem_write_data_reg_29),
	.prn(vcc));
defparam \mem_write_data_reg[29] .is_wysiwyg = "true";
defparam \mem_write_data_reg[29] .power_up = "low";

dffeas \mem_write_data_reg[28] (
	.clk(clk_clk),
	.d(avl_mem_writedata_28),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(mem_write_data_reg_28),
	.prn(vcc));
defparam \mem_write_data_reg[28] .is_wysiwyg = "true";
defparam \mem_write_data_reg[28] .power_up = "low";

dffeas \mem_write_data_reg[27] (
	.clk(clk_clk),
	.d(avl_mem_writedata_27),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(mem_write_data_reg_27),
	.prn(vcc));
defparam \mem_write_data_reg[27] .is_wysiwyg = "true";
defparam \mem_write_data_reg[27] .power_up = "low";

cycloneive_lcell_comb \cmd_data[11] (
	.dataa(\mem_write_data_reg[11]~q ),
	.datab(\cmd_data[11]~4_combout ),
	.datac(\cmd_data[8]~88_combout ),
	.datad(\cmd_data[11]~7_combout ),
	.cin(gnd),
	.combout(cmd_data_11),
	.cout());
defparam \cmd_data[11] .lut_mask = 16'hCFA0;
defparam \cmd_data[11] .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~1 (
	.dataa(mem_byteenable_reg_0),
	.datab(mem_byteenable_reg_3),
	.datac(mem_byteenable_reg_2),
	.datad(mem_byteenable_reg_1),
	.cin(gnd),
	.combout(Add1),
	.cout());
defparam \Add1~1 .lut_mask = 16'h6996;
defparam \Add1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector20~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(current_stateSTATE_WR_CMD),
	.datad(current_stateSTATE_READ_CMD),
	.cin(gnd),
	.combout(Selector20),
	.cout());
defparam \Selector20~0 .lut_mask = 16'h000F;
defparam \Selector20~0 .sum_lutc_input = "datac";

dffeas \mem_write_data_reg[18] (
	.clk(clk_clk),
	.d(avl_mem_writedata_18),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(mem_write_data_reg_18),
	.prn(vcc));
defparam \mem_write_data_reg[18] .is_wysiwyg = "true";
defparam \mem_write_data_reg[18] .power_up = "low";

cycloneive_lcell_comb \Add1~2 (
	.dataa(mem_byteenable_reg_0),
	.datab(mem_byteenable_reg_3),
	.datac(mem_byteenable_reg_2),
	.datad(mem_byteenable_reg_1),
	.cin(gnd),
	.combout(Add11),
	.cout());
defparam \Add1~2 .lut_mask = 16'h7EE8;
defparam \Add1~2 .sum_lutc_input = "datac";

dffeas \mem_write_data_reg[19] (
	.clk(clk_clk),
	.d(avl_mem_writedata_19),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(mem_write_data_reg_19),
	.prn(vcc));
defparam \mem_write_data_reg[19] .is_wysiwyg = "true";
defparam \mem_write_data_reg[19] .power_up = "low";

dffeas \mem_write_data_reg[21] (
	.clk(clk_clk),
	.d(avl_mem_writedata_21),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(mem_write_data_reg_21),
	.prn(vcc));
defparam \mem_write_data_reg[21] .is_wysiwyg = "true";
defparam \mem_write_data_reg[21] .power_up = "low";

dffeas \mem_burstcount_reg[1] (
	.clk(clk_clk),
	.d(mem_burstcount[1]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_burstcount_reg_1),
	.prn(vcc));
defparam \mem_burstcount_reg[1] .is_wysiwyg = "true";
defparam \mem_burstcount_reg[1] .power_up = "low";

dffeas \mem_write_data_reg[20] (
	.clk(clk_clk),
	.d(avl_mem_writedata_20),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(mem_write_data_reg_20),
	.prn(vcc));
defparam \mem_write_data_reg[20] .is_wysiwyg = "true";
defparam \mem_write_data_reg[20] .power_up = "low";

dffeas \mem_burstcount_reg[0] (
	.clk(clk_clk),
	.d(mem_burstcount[0]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_burstcount_reg_0),
	.prn(vcc));
defparam \mem_burstcount_reg[0] .is_wysiwyg = "true";
defparam \mem_burstcount_reg[0] .power_up = "low";

dffeas \mem_write_data_reg[22] (
	.clk(clk_clk),
	.d(avl_mem_writedata_22),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(mem_write_data_reg_22),
	.prn(vcc));
defparam \mem_write_data_reg[22] .is_wysiwyg = "true";
defparam \mem_write_data_reg[22] .power_up = "low";

dffeas \mem_burstcount_reg[2] (
	.clk(clk_clk),
	.d(mem_burstcount[2]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_burstcount_reg_2),
	.prn(vcc));
defparam \mem_burstcount_reg[2] .is_wysiwyg = "true";
defparam \mem_burstcount_reg[2] .power_up = "low";

dffeas \mem_write_data_reg[23] (
	.clk(clk_clk),
	.d(avl_mem_writedata_23),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(mem_write_data_reg_23),
	.prn(vcc));
defparam \mem_write_data_reg[23] .is_wysiwyg = "true";
defparam \mem_write_data_reg[23] .power_up = "low";

dffeas \mem_burstcount_reg[3] (
	.clk(clk_clk),
	.d(mem_burstcount[3]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_burstcount_reg_3),
	.prn(vcc));
defparam \mem_burstcount_reg[3] .is_wysiwyg = "true";
defparam \mem_burstcount_reg[3] .power_up = "low";

dffeas \mem_write_data_reg[24] (
	.clk(clk_clk),
	.d(avl_mem_writedata_24),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(mem_write_data_reg_24),
	.prn(vcc));
defparam \mem_write_data_reg[24] .is_wysiwyg = "true";
defparam \mem_write_data_reg[24] .power_up = "low";

dffeas \mem_burstcount_reg[4] (
	.clk(clk_clk),
	.d(mem_burstcount[4]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_burstcount_reg_4),
	.prn(vcc));
defparam \mem_burstcount_reg[4] .is_wysiwyg = "true";
defparam \mem_burstcount_reg[4] .power_up = "low";

dffeas \mem_write_data_reg[25] (
	.clk(clk_clk),
	.d(avl_mem_writedata_25),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(mem_write_data_reg_25),
	.prn(vcc));
defparam \mem_write_data_reg[25] .is_wysiwyg = "true";
defparam \mem_write_data_reg[25] .power_up = "low";

dffeas \mem_burstcount_reg[5] (
	.clk(clk_clk),
	.d(mem_burstcount[5]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_burstcount_reg_5),
	.prn(vcc));
defparam \mem_burstcount_reg[5] .is_wysiwyg = "true";
defparam \mem_burstcount_reg[5] .power_up = "low";

dffeas \mem_write_data_reg[26] (
	.clk(clk_clk),
	.d(avl_mem_writedata_26),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(mem_write_data_reg_26),
	.prn(vcc));
defparam \mem_write_data_reg[26] .is_wysiwyg = "true";
defparam \mem_write_data_reg[26] .power_up = "low";

dffeas \mem_burstcount_reg[6] (
	.clk(clk_clk),
	.d(mem_burstcount[6]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_burstcount_reg_6),
	.prn(vcc));
defparam \mem_burstcount_reg[6] .is_wysiwyg = "true";
defparam \mem_burstcount_reg[6] .power_up = "low";

cycloneive_lcell_comb \cmd_data[10] (
	.dataa(\mem_write_data_reg[10]~q ),
	.datab(\cmd_data[10]~8_combout ),
	.datac(\cmd_data[8]~88_combout ),
	.datad(\cmd_data[10]~9_combout ),
	.cin(gnd),
	.combout(cmd_data_10),
	.cout());
defparam \cmd_data[10] .lut_mask = 16'hCFA0;
defparam \cmd_data[10] .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[8] (
	.dataa(\mem_write_data_reg[8]~q ),
	.datab(\cmd_data[8]~10_combout ),
	.datac(\cmd_data[8]~88_combout ),
	.datad(\cmd_data[8]~11_combout ),
	.cin(gnd),
	.combout(cmd_data_8),
	.cout());
defparam \cmd_data[8] .lut_mask = 16'hCFA0;
defparam \cmd_data[8] .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[13] (
	.dataa(\mem_write_data_reg[13]~q ),
	.datab(\cmd_data[13]~12_combout ),
	.datac(\cmd_data[8]~88_combout ),
	.datad(\cmd_data[13]~13_combout ),
	.cin(gnd),
	.combout(cmd_data_13),
	.cout());
defparam \cmd_data[13] .lut_mask = 16'hCFA0;
defparam \cmd_data[13] .sum_lutc_input = "datac";

dffeas \mem_write_data_reg[17] (
	.clk(clk_clk),
	.d(avl_mem_writedata_17),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(mem_write_data_reg_17),
	.prn(vcc));
defparam \mem_write_data_reg[17] .is_wysiwyg = "true";
defparam \mem_write_data_reg[17] .power_up = "low";

dffeas \mem_write_data_reg[16] (
	.clk(clk_clk),
	.d(avl_mem_writedata_16),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(mem_write_data_reg_16),
	.prn(vcc));
defparam \mem_write_data_reg[16] .is_wysiwyg = "true";
defparam \mem_write_data_reg[16] .power_up = "low";

dffeas \mem_write_data_reg[31] (
	.clk(clk_clk),
	.d(avl_mem_writedata_31),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(mem_write_data_reg_31),
	.prn(vcc));
defparam \mem_write_data_reg[31] .is_wysiwyg = "true";
defparam \mem_write_data_reg[31] .power_up = "low";

cycloneive_lcell_comb \cmd_data[15] (
	.dataa(\mem_write_data_reg[15]~q ),
	.datab(\cmd_data[15]~14_combout ),
	.datac(\cmd_data[14]~89_combout ),
	.datad(\cmd_data[15]~17_combout ),
	.cin(gnd),
	.combout(cmd_data_15),
	.cout());
defparam \cmd_data[15] .lut_mask = 16'hCFA0;
defparam \cmd_data[15] .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[14] (
	.dataa(\mem_write_data_reg[14]~q ),
	.datab(\cmd_data[14]~18_combout ),
	.datac(\cmd_data[14]~89_combout ),
	.datad(\cmd_data[14]~20_combout ),
	.cin(gnd),
	.combout(cmd_data_14),
	.cout());
defparam \cmd_data[14] .lut_mask = 16'hCFA0;
defparam \cmd_data[14] .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[9] (
	.dataa(\mem_write_data_reg[9]~q ),
	.datab(\cmd_data[9]~21_combout ),
	.datac(\cmd_data[8]~88_combout ),
	.datad(\cmd_data[9]~22_combout ),
	.cin(gnd),
	.combout(cmd_data_9),
	.cout());
defparam \cmd_data[9] .lut_mask = 16'hCFA0;
defparam \cmd_data[9] .sum_lutc_input = "datac";

dffeas \mem_addr_reg[6] (
	.clk(clk_clk),
	.d(mem_addr[6]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_addr_reg_6),
	.prn(vcc));
defparam \mem_addr_reg[6] .is_wysiwyg = "true";
defparam \mem_addr_reg[6] .power_up = "low";

dffeas \mem_addr_reg[14] (
	.clk(clk_clk),
	.d(mem_addr[14]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_addr_reg_14),
	.prn(vcc));
defparam \mem_addr_reg[14] .is_wysiwyg = "true";
defparam \mem_addr_reg[14] .power_up = "low";

cycloneive_lcell_comb \addr_bytes_xip[0]~0 (
	.dataa(mem_byteenable_reg_0),
	.datab(mem_byteenable_reg_1),
	.datac(mem_byteenable_reg_2),
	.datad(mem_byteenable_reg_3),
	.cin(gnd),
	.combout(addr_bytes_xip_0),
	.cout());
defparam \addr_bytes_xip[0]~0 .lut_mask = 16'h0104;
defparam \addr_bytes_xip[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[0]~36 (
	.dataa(\cmd_data[0]~23_combout ),
	.datab(csr_wr_inst_data_8),
	.datac(\cmd_data[2]~24_combout ),
	.datad(\cmd_data[0]~35_combout ),
	.cin(gnd),
	.combout(cmd_data_0),
	.cout());
defparam \cmd_data[0]~36 .lut_mask = 16'hFC0A;
defparam \cmd_data[0]~36 .sum_lutc_input = "datac";

dffeas \mem_addr_reg[10] (
	.clk(clk_clk),
	.d(mem_addr[10]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_addr_reg_10),
	.prn(vcc));
defparam \mem_addr_reg[10] .is_wysiwyg = "true";
defparam \mem_addr_reg[10] .power_up = "low";

dffeas \mem_addr_reg[18] (
	.clk(clk_clk),
	.d(mem_addr[18]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_addr_reg_18),
	.prn(vcc));
defparam \mem_addr_reg[18] .is_wysiwyg = "true";
defparam \mem_addr_reg[18] .power_up = "low";

dffeas \mem_addr_reg[2] (
	.clk(clk_clk),
	.d(mem_addr[2]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_addr_reg_2),
	.prn(vcc));
defparam \mem_addr_reg[2] .is_wysiwyg = "true";
defparam \mem_addr_reg[2] .power_up = "low";

cycloneive_lcell_comb \cmd_data[4]~43 (
	.dataa(\cmd_data[4]~37_combout ),
	.datab(csr_wr_inst_data_12),
	.datac(\cmd_data[2]~24_combout ),
	.datad(\cmd_data[4]~42_combout ),
	.cin(gnd),
	.combout(cmd_data_4),
	.cout());
defparam \cmd_data[4]~43 .lut_mask = 16'hF30A;
defparam \cmd_data[4]~43 .sum_lutc_input = "datac";

dffeas \mem_addr_reg[8] (
	.clk(clk_clk),
	.d(mem_addr[8]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_addr_reg_8),
	.prn(vcc));
defparam \mem_addr_reg[8] .is_wysiwyg = "true";
defparam \mem_addr_reg[8] .power_up = "low";

dffeas \mem_addr_reg[16] (
	.clk(clk_clk),
	.d(mem_addr[16]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_addr_reg_16),
	.prn(vcc));
defparam \mem_addr_reg[16] .is_wysiwyg = "true";
defparam \mem_addr_reg[16] .power_up = "low";

dffeas \mem_addr_reg[0] (
	.clk(clk_clk),
	.d(mem_addr[0]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_addr_reg_0),
	.prn(vcc));
defparam \mem_addr_reg[0] .is_wysiwyg = "true";
defparam \mem_addr_reg[0] .power_up = "low";

cycloneive_lcell_comb \cmd_data[2]~50 (
	.dataa(\cmd_data[2]~44_combout ),
	.datab(csr_wr_inst_data_10),
	.datac(\cmd_data[2]~24_combout ),
	.datad(\cmd_data[2]~49_combout ),
	.cin(gnd),
	.combout(cmd_data_2),
	.cout());
defparam \cmd_data[2]~50 .lut_mask = 16'hFC0A;
defparam \cmd_data[2]~50 .sum_lutc_input = "datac";

dffeas \mem_addr_reg[15] (
	.clk(clk_clk),
	.d(mem_addr[15]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_addr_reg_15),
	.prn(vcc));
defparam \mem_addr_reg[15] .is_wysiwyg = "true";
defparam \mem_addr_reg[15] .power_up = "low";

dffeas \mem_addr_reg[7] (
	.clk(clk_clk),
	.d(mem_addr[7]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_addr_reg_7),
	.prn(vcc));
defparam \mem_addr_reg[7] .is_wysiwyg = "true";
defparam \mem_addr_reg[7] .power_up = "low";

cycloneive_lcell_comb \WideOr19~0 (
	.dataa(mem_byteenable_reg_0),
	.datab(mem_byteenable_reg_1),
	.datac(mem_byteenable_reg_2),
	.datad(mem_byteenable_reg_3),
	.cin(gnd),
	.combout(WideOr19),
	.cout());
defparam \WideOr19~0 .lut_mask = 16'h1110;
defparam \WideOr19~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[1]~57 (
	.dataa(\cmd_data[1]~51_combout ),
	.datab(csr_wr_inst_data_9),
	.datac(\cmd_data[2]~24_combout ),
	.datad(\cmd_data[1]~56_combout ),
	.cin(gnd),
	.combout(cmd_data_1),
	.cout());
defparam \cmd_data[1]~57 .lut_mask = 16'hFC0A;
defparam \cmd_data[1]~57 .sum_lutc_input = "datac";

dffeas \mem_addr_reg[17] (
	.clk(clk_clk),
	.d(mem_addr[17]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_addr_reg_17),
	.prn(vcc));
defparam \mem_addr_reg[17] .is_wysiwyg = "true";
defparam \mem_addr_reg[17] .power_up = "low";

dffeas \mem_addr_reg[9] (
	.clk(clk_clk),
	.d(mem_addr[9]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_addr_reg_9),
	.prn(vcc));
defparam \mem_addr_reg[9] .is_wysiwyg = "true";
defparam \mem_addr_reg[9] .power_up = "low";

dffeas \mem_addr_reg[1] (
	.clk(clk_clk),
	.d(mem_addr[1]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_addr_reg_1),
	.prn(vcc));
defparam \mem_addr_reg[1] .is_wysiwyg = "true";
defparam \mem_addr_reg[1] .power_up = "low";

cycloneive_lcell_comb \cmd_data[3]~64 (
	.dataa(\cmd_data[3]~58_combout ),
	.datab(csr_wr_inst_data_11),
	.datac(\cmd_data[2]~24_combout ),
	.datad(\cmd_data[3]~63_combout ),
	.cin(gnd),
	.combout(cmd_data_3),
	.cout());
defparam \cmd_data[3]~64 .lut_mask = 16'hFC0A;
defparam \cmd_data[3]~64 .sum_lutc_input = "datac";

dffeas \mem_addr_reg[19] (
	.clk(clk_clk),
	.d(mem_addr[19]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_addr_reg_19),
	.prn(vcc));
defparam \mem_addr_reg[19] .is_wysiwyg = "true";
defparam \mem_addr_reg[19] .power_up = "low";

dffeas \mem_addr_reg[11] (
	.clk(clk_clk),
	.d(mem_addr[11]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_addr_reg_11),
	.prn(vcc));
defparam \mem_addr_reg[11] .is_wysiwyg = "true";
defparam \mem_addr_reg[11] .power_up = "low";

dffeas \mem_addr_reg[3] (
	.clk(clk_clk),
	.d(mem_addr[3]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_addr_reg_3),
	.prn(vcc));
defparam \mem_addr_reg[3] .is_wysiwyg = "true";
defparam \mem_addr_reg[3] .power_up = "low";

cycloneive_lcell_comb \cmd_data[5]~71 (
	.dataa(\cmd_data[5]~65_combout ),
	.datab(csr_wr_inst_data_13),
	.datac(\cmd_data[2]~24_combout ),
	.datad(\cmd_data[5]~70_combout ),
	.cin(gnd),
	.combout(cmd_data_5),
	.cout());
defparam \cmd_data[5]~71 .lut_mask = 16'hF30A;
defparam \cmd_data[5]~71 .sum_lutc_input = "datac";

dffeas \mem_addr_reg[12] (
	.clk(clk_clk),
	.d(mem_addr[12]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_addr_reg_12),
	.prn(vcc));
defparam \mem_addr_reg[12] .is_wysiwyg = "true";
defparam \mem_addr_reg[12] .power_up = "low";

dffeas \mem_addr_reg[20] (
	.clk(clk_clk),
	.d(mem_addr[20]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_addr_reg_20),
	.prn(vcc));
defparam \mem_addr_reg[20] .is_wysiwyg = "true";
defparam \mem_addr_reg[20] .power_up = "low";

dffeas \mem_addr_reg[4] (
	.clk(clk_clk),
	.d(mem_addr[4]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_addr_reg_4),
	.prn(vcc));
defparam \mem_addr_reg[4] .is_wysiwyg = "true";
defparam \mem_addr_reg[4] .power_up = "low";

cycloneive_lcell_comb \cmd_data[6]~78 (
	.dataa(\cmd_data[6]~72_combout ),
	.datab(csr_wr_inst_data_14),
	.datac(\cmd_data[2]~24_combout ),
	.datad(\cmd_data[6]~77_combout ),
	.cin(gnd),
	.combout(cmd_data_6),
	.cout());
defparam \cmd_data[6]~78 .lut_mask = 16'hF30A;
defparam \cmd_data[6]~78 .sum_lutc_input = "datac";

dffeas \mem_addr_reg[13] (
	.clk(clk_clk),
	.d(mem_addr[13]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_addr_reg_13),
	.prn(vcc));
defparam \mem_addr_reg[13] .is_wysiwyg = "true";
defparam \mem_addr_reg[13] .power_up = "low";

dffeas \mem_addr_reg[5] (
	.clk(clk_clk),
	.d(mem_addr[5]),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_byteenable_reg[0]~3_combout ),
	.q(mem_addr_reg_5),
	.prn(vcc));
defparam \mem_addr_reg[5] .is_wysiwyg = "true";
defparam \mem_addr_reg[5] .power_up = "low";

cycloneive_lcell_comb \cmd_data[7]~85 (
	.dataa(\cmd_data[7]~79_combout ),
	.datab(csr_wr_inst_data_15),
	.datac(\cmd_data[2]~24_combout ),
	.datad(\cmd_data[7]~84_combout ),
	.cin(gnd),
	.combout(cmd_data_7),
	.cout());
defparam \cmd_data[7]~85 .lut_mask = 16'hFC0A;
defparam \cmd_data[7]~85 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[12] (
	.dataa(\mem_write_data_reg[12]~q ),
	.datab(\cmd_data[12]~86_combout ),
	.datac(\cmd_data[8]~88_combout ),
	.datad(\cmd_data[12]~87_combout ),
	.cin(gnd),
	.combout(cmd_data_12),
	.cout());
defparam \cmd_data[12] .lut_mask = 16'hCFA0;
defparam \cmd_data[12] .sum_lutc_input = "datac";

cycloneive_lcell_comb \always0~0 (
	.dataa(in_cmd_channel_reg_0),
	.datab(stateST_SEND_DUMMY_RSP),
	.datac(out_valid),
	.datad(out_endofpacket),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
defparam \always0~0 .lut_mask = 16'hA888;
defparam \always0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector8~0 (
	.dataa(current_stateSTATE_POLL_CMD),
	.datab(sink0_ready),
	.datac(\current_state.STATE_POLL_RSP~q ),
	.datad(\always0~0_combout ),
	.cin(gnd),
	.combout(\Selector8~0_combout ),
	.cout());
defparam \Selector8~0 .lut_mask = 16'h88F8;
defparam \Selector8~0 .sum_lutc_input = "datac";

dffeas \current_state.STATE_POLL_RSP (
	.clk(clk_clk),
	.d(\Selector8~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\current_state.STATE_POLL_RSP~q ),
	.prn(vcc));
defparam \current_state.STATE_POLL_RSP .is_wysiwyg = "true";
defparam \current_state.STATE_POLL_RSP .power_up = "low";

cycloneive_lcell_comb \Equal3~0 (
	.dataa(csr_wr_inst_data_12),
	.datab(csr_wr_inst_data_13),
	.datac(csr_wr_inst_data_14),
	.datad(csr_wr_inst_data_15),
	.cin(gnd),
	.combout(\Equal3~0_combout ),
	.cout());
defparam \Equal3~0 .lut_mask = 16'h0001;
defparam \Equal3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal3~1 (
	.dataa(csr_wr_inst_data_8),
	.datab(csr_wr_inst_data_9),
	.datac(csr_wr_inst_data_10),
	.datad(csr_wr_inst_data_11),
	.cin(gnd),
	.combout(\Equal3~1_combout ),
	.cout());
defparam \Equal3~1 .lut_mask = 16'h0001;
defparam \Equal3~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \busy~0 (
	.dataa(out_rsp_data_7),
	.datab(out_rsp_data_0),
	.datac(\Equal3~0_combout ),
	.datad(\Equal3~1_combout ),
	.cin(gnd),
	.combout(\busy~0_combout ),
	.cout());
defparam \busy~0 .lut_mask = 16'h5CCC;
defparam \busy~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector12~0 (
	.dataa(\always0~0_combout ),
	.datab(current_stateSTATE_READ_DATA),
	.datac(\current_state.STATE_POLL_RSP~q ),
	.datad(\busy~0_combout ),
	.cin(gnd),
	.combout(\Selector12~0_combout ),
	.cout());
defparam \Selector12~0 .lut_mask = 16'h88A8;
defparam \Selector12~0 .sum_lutc_input = "datac";

dffeas \current_state.STATE_COMPLETE (
	.clk(clk_clk),
	.d(\Selector12~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\current_state.STATE_COMPLETE~q ),
	.prn(vcc));
defparam \current_state.STATE_COMPLETE .is_wysiwyg = "true";
defparam \current_state.STATE_COMPLETE .power_up = "low";

cycloneive_lcell_comb \burstcount_register[0]~7 (
	.dataa(\internal_burstcount[0]~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\burstcount_register[0]~7_combout ),
	.cout(\burstcount_register[0]~8 ));
defparam \burstcount_register[0]~7 .lut_mask = 16'h55AA;
defparam \burstcount_register[0]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(avl_mem_byteenable_0),
	.datab(avl_mem_byteenable_1),
	.datac(avl_mem_byteenable_2),
	.datad(avl_mem_byteenable_3),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h0001;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \sop_enable~0 (
	.dataa(\Equal2~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\sop_enable~0_combout ),
	.cout());
defparam \sop_enable~0 .lut_mask = 16'h5555;
defparam \sop_enable~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_wr_combi~0 (
	.dataa(hold_waitrequest1),
	.datab(avl_mem_write),
	.datac(\current_state.STATE_IDLE~q ),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\mem_wr_combi~0_combout ),
	.cout());
defparam \mem_wr_combi~0 .lut_mask = 16'h0008;
defparam \mem_wr_combi~0 .sum_lutc_input = "datac";

dffeas sop_enable(
	.clk(clk_clk),
	.d(\sop_enable~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(\sop_enable~q ),
	.prn(vcc));
defparam sop_enable.is_wysiwyg = "true";
defparam sop_enable.power_up = "low";

cycloneive_lcell_comb \burstcount_register~9 (
	.dataa(mem_waitrequest),
	.datab(avl_mem_write),
	.datac(\Equal0~0_combout ),
	.datad(\sop_enable~q ),
	.cin(gnd),
	.combout(\burstcount_register~9_combout ),
	.cout());
defparam \burstcount_register~9 .lut_mask = 16'h08FF;
defparam \burstcount_register~9 .sum_lutc_input = "datac";

dffeas \burstcount_register[0] (
	.clk(clk_clk),
	.d(\burstcount_register[0]~7_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\burstcount_register~9_combout ),
	.q(\burstcount_register[0]~q ),
	.prn(vcc));
defparam \burstcount_register[0] .is_wysiwyg = "true";
defparam \burstcount_register[0] .power_up = "low";

cycloneive_lcell_comb \internal_burstcount[0]~0 (
	.dataa(\burstcount_register[0]~q ),
	.datab(mem_burstcount[0]),
	.datac(gnd),
	.datad(\sop_enable~q ),
	.cin(gnd),
	.combout(\internal_burstcount[0]~0_combout ),
	.cout());
defparam \internal_burstcount[0]~0 .lut_mask = 16'hAACC;
defparam \internal_burstcount[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \burstcount_register[1]~10 (
	.dataa(\internal_burstcount[1]~3_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\burstcount_register[0]~8 ),
	.combout(\burstcount_register[1]~10_combout ),
	.cout(\burstcount_register[1]~11 ));
defparam \burstcount_register[1]~10 .lut_mask = 16'hA505;
defparam \burstcount_register[1]~10 .sum_lutc_input = "cin";

dffeas \burstcount_register[1] (
	.clk(clk_clk),
	.d(\burstcount_register[1]~10_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\burstcount_register~9_combout ),
	.q(\burstcount_register[1]~q ),
	.prn(vcc));
defparam \burstcount_register[1] .is_wysiwyg = "true";
defparam \burstcount_register[1] .power_up = "low";

cycloneive_lcell_comb \internal_burstcount[1]~3 (
	.dataa(\burstcount_register[1]~q ),
	.datab(mem_burstcount[1]),
	.datac(gnd),
	.datad(\sop_enable~q ),
	.cin(gnd),
	.combout(\internal_burstcount[1]~3_combout ),
	.cout());
defparam \internal_burstcount[1]~3 .lut_mask = 16'hAACC;
defparam \internal_burstcount[1]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \burstcount_register[2]~12 (
	.dataa(\internal_burstcount[2]~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\burstcount_register[1]~11 ),
	.combout(\burstcount_register[2]~12_combout ),
	.cout(\burstcount_register[2]~13 ));
defparam \burstcount_register[2]~12 .lut_mask = 16'h5AAF;
defparam \burstcount_register[2]~12 .sum_lutc_input = "cin";

dffeas \burstcount_register[2] (
	.clk(clk_clk),
	.d(\burstcount_register[2]~12_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\burstcount_register~9_combout ),
	.q(\burstcount_register[2]~q ),
	.prn(vcc));
defparam \burstcount_register[2] .is_wysiwyg = "true";
defparam \burstcount_register[2] .power_up = "low";

cycloneive_lcell_comb \internal_burstcount[2]~2 (
	.dataa(\burstcount_register[2]~q ),
	.datab(mem_burstcount[2]),
	.datac(gnd),
	.datad(\sop_enable~q ),
	.cin(gnd),
	.combout(\internal_burstcount[2]~2_combout ),
	.cout());
defparam \internal_burstcount[2]~2 .lut_mask = 16'hAACC;
defparam \internal_burstcount[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \burstcount_register[3]~14 (
	.dataa(\internal_burstcount[3]~6_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\burstcount_register[2]~13 ),
	.combout(\burstcount_register[3]~14_combout ),
	.cout(\burstcount_register[3]~15 ));
defparam \burstcount_register[3]~14 .lut_mask = 16'hA505;
defparam \burstcount_register[3]~14 .sum_lutc_input = "cin";

dffeas \burstcount_register[3] (
	.clk(clk_clk),
	.d(\burstcount_register[3]~14_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\burstcount_register~9_combout ),
	.q(\burstcount_register[3]~q ),
	.prn(vcc));
defparam \burstcount_register[3] .is_wysiwyg = "true";
defparam \burstcount_register[3] .power_up = "low";

cycloneive_lcell_comb \internal_burstcount[3]~6 (
	.dataa(\burstcount_register[3]~q ),
	.datab(mem_burstcount[3]),
	.datac(gnd),
	.datad(\sop_enable~q ),
	.cin(gnd),
	.combout(\internal_burstcount[3]~6_combout ),
	.cout());
defparam \internal_burstcount[3]~6 .lut_mask = 16'hAACC;
defparam \internal_burstcount[3]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \burstcount_register[4]~16 (
	.dataa(\internal_burstcount[4]~5_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\burstcount_register[3]~15 ),
	.combout(\burstcount_register[4]~16_combout ),
	.cout(\burstcount_register[4]~17 ));
defparam \burstcount_register[4]~16 .lut_mask = 16'h5AAF;
defparam \burstcount_register[4]~16 .sum_lutc_input = "cin";

dffeas \burstcount_register[4] (
	.clk(clk_clk),
	.d(\burstcount_register[4]~16_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\burstcount_register~9_combout ),
	.q(\burstcount_register[4]~q ),
	.prn(vcc));
defparam \burstcount_register[4] .is_wysiwyg = "true";
defparam \burstcount_register[4] .power_up = "low";

cycloneive_lcell_comb \internal_burstcount[4]~5 (
	.dataa(\burstcount_register[4]~q ),
	.datab(mem_burstcount[4]),
	.datac(gnd),
	.datad(\sop_enable~q ),
	.cin(gnd),
	.combout(\internal_burstcount[4]~5_combout ),
	.cout());
defparam \internal_burstcount[4]~5 .lut_mask = 16'hAACC;
defparam \internal_burstcount[4]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \burstcount_register[5]~18 (
	.dataa(\internal_burstcount[5]~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\burstcount_register[4]~17 ),
	.combout(\burstcount_register[5]~18_combout ),
	.cout(\burstcount_register[5]~19 ));
defparam \burstcount_register[5]~18 .lut_mask = 16'hA505;
defparam \burstcount_register[5]~18 .sum_lutc_input = "cin";

dffeas \burstcount_register[5] (
	.clk(clk_clk),
	.d(\burstcount_register[5]~18_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\burstcount_register~9_combout ),
	.q(\burstcount_register[5]~q ),
	.prn(vcc));
defparam \burstcount_register[5] .is_wysiwyg = "true";
defparam \burstcount_register[5] .power_up = "low";

cycloneive_lcell_comb \internal_burstcount[5]~4 (
	.dataa(\burstcount_register[5]~q ),
	.datab(mem_burstcount[5]),
	.datac(gnd),
	.datad(\sop_enable~q ),
	.cin(gnd),
	.combout(\internal_burstcount[5]~4_combout ),
	.cout());
defparam \internal_burstcount[5]~4 .lut_mask = 16'hAACC;
defparam \internal_burstcount[5]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \burstcount_register[6]~20 (
	.dataa(\internal_burstcount[6]~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\burstcount_register[5]~19 ),
	.combout(\burstcount_register[6]~20_combout ),
	.cout());
defparam \burstcount_register[6]~20 .lut_mask = 16'h5A5A;
defparam \burstcount_register[6]~20 .sum_lutc_input = "cin";

dffeas \burstcount_register[6] (
	.clk(clk_clk),
	.d(\burstcount_register[6]~20_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\burstcount_register~9_combout ),
	.q(\burstcount_register[6]~q ),
	.prn(vcc));
defparam \burstcount_register[6] .is_wysiwyg = "true";
defparam \burstcount_register[6] .power_up = "low";

cycloneive_lcell_comb \internal_burstcount[6]~1 (
	.dataa(\burstcount_register[6]~q ),
	.datab(mem_burstcount[6]),
	.datac(gnd),
	.datad(\sop_enable~q ),
	.cin(gnd),
	.combout(\internal_burstcount[6]~1_combout ),
	.cout());
defparam \internal_burstcount[6]~1 .lut_mask = 16'hAACC;
defparam \internal_burstcount[6]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal2~0 (
	.dataa(\internal_burstcount[0]~0_combout ),
	.datab(\internal_burstcount[6]~1_combout ),
	.datac(\internal_burstcount[2]~2_combout ),
	.datad(\internal_burstcount[1]~3_combout ),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
defparam \Equal2~0 .lut_mask = 16'h0002;
defparam \Equal2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal2~1 (
	.dataa(\Equal2~0_combout ),
	.datab(\internal_burstcount[5]~4_combout ),
	.datac(\internal_burstcount[4]~5_combout ),
	.datad(\internal_burstcount[3]~6_combout ),
	.cin(gnd),
	.combout(\Equal2~1_combout ),
	.cout());
defparam \Equal2~1 .lut_mask = 16'h0002;
defparam \Equal2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector0~0 (
	.dataa(avl_mem_write),
	.datab(gnd),
	.datac(\avst_fifo_inst|avst_fifo|full~q ),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
defparam \Selector0~0 .lut_mask = 16'h000A;
defparam \Selector0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector0~1 (
	.dataa(hold_waitrequest1),
	.datab(avl_mem_read),
	.datac(\Equal2~1_combout ),
	.datad(\Selector0~0_combout ),
	.cin(gnd),
	.combout(\Selector0~1_combout ),
	.cout());
defparam \Selector0~1 .lut_mask = 16'hA888;
defparam \Selector0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector0~2 (
	.dataa(\current_state.STATE_COMPLETE~q ),
	.datab(gnd),
	.datac(\current_state.STATE_IDLE~q ),
	.datad(\Selector0~1_combout ),
	.cin(gnd),
	.combout(\Selector0~2_combout ),
	.cout());
defparam \Selector0~2 .lut_mask = 16'h5550;
defparam \Selector0~2 .sum_lutc_input = "datac";

dffeas \current_state.STATE_IDLE (
	.clk(clk_clk),
	.d(\Selector0~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\current_state.STATE_IDLE~q ),
	.prn(vcc));
defparam \current_state.STATE_IDLE .is_wysiwyg = "true";
defparam \current_state.STATE_IDLE .power_up = "low";

cycloneive_lcell_comb \mem_rddatavalid~0 (
	.dataa(current_stateSTATE_READ_DATA),
	.datab(in_cmd_channel_reg_0),
	.datac(out_valid),
	.datad(stateST_SEND_DUMMY_RSP),
	.cin(gnd),
	.combout(\mem_rddatavalid~0_combout ),
	.cout());
defparam \mem_rddatavalid~0 .lut_mask = 16'h8880;
defparam \mem_rddatavalid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector11~0 (
	.dataa(current_stateSTATE_READ_CMD),
	.datab(sink0_ready),
	.datac(current_stateSTATE_READ_DATA),
	.datad(\always0~0_combout ),
	.cin(gnd),
	.combout(\Selector11~0_combout ),
	.cout());
defparam \Selector11~0 .lut_mask = 16'h88F8;
defparam \Selector11~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~0 (
	.dataa(current_stateSTATE_STATUS_CMD),
	.datab(sink0_ready),
	.datac(\current_state.STATE_STATUS_RSP~q ),
	.datad(\always0~0_combout ),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
defparam \Selector2~0 .lut_mask = 16'h88F8;
defparam \Selector2~0 .sum_lutc_input = "datac";

dffeas \current_state.STATE_STATUS_RSP (
	.clk(clk_clk),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\current_state.STATE_STATUS_RSP~q ),
	.prn(vcc));
defparam \current_state.STATE_STATUS_RSP .is_wysiwyg = "true";
defparam \current_state.STATE_STATUS_RSP .power_up = "low";

cycloneive_lcell_comb \Selector3~0 (
	.dataa(\current_state.STATE_STATUS_RSP~q ),
	.datab(gnd),
	.datac(out_valid),
	.datad(out_data_0),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
defparam \Selector3~0 .lut_mask = 16'h0AAA;
defparam \Selector3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector3~1 (
	.dataa(\always0~0_combout ),
	.datab(\Selector3~0_combout ),
	.datac(\current_state.STATE_WRENABLE_CMD~q ),
	.datad(sink0_ready),
	.cin(gnd),
	.combout(\Selector3~1_combout ),
	.cout());
defparam \Selector3~1 .lut_mask = 16'h88F8;
defparam \Selector3~1 .sum_lutc_input = "datac";

dffeas \current_state.STATE_WRENABLE_CMD (
	.clk(clk_clk),
	.d(\Selector3~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\current_state.STATE_WRENABLE_CMD~q ),
	.prn(vcc));
defparam \current_state.STATE_WRENABLE_CMD .is_wysiwyg = "true";
defparam \current_state.STATE_WRENABLE_CMD .power_up = "low";

cycloneive_lcell_comb \Selector4~0 (
	.dataa(\current_state.STATE_WRENABLE_CMD~q ),
	.datab(sink0_ready),
	.datac(\current_state.STATE_WRENABLE_RSP~q ),
	.datad(\always0~0_combout ),
	.cin(gnd),
	.combout(\Selector4~0_combout ),
	.cout());
defparam \Selector4~0 .lut_mask = 16'h88F8;
defparam \Selector4~0 .sum_lutc_input = "datac";

dffeas \current_state.STATE_WRENABLE_RSP (
	.clk(clk_clk),
	.d(\Selector4~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\current_state.STATE_WRENABLE_RSP~q ),
	.prn(vcc));
defparam \current_state.STATE_WRENABLE_RSP .is_wysiwyg = "true";
defparam \current_state.STATE_WRENABLE_RSP .power_up = "low";

cycloneive_lcell_comb \Selector5~0 (
	.dataa(\always0~0_combout ),
	.datab(\current_state.STATE_WRENABLE_RSP~q ),
	.datac(current_stateSTATE_WR_CMD),
	.datad(sink0_ready),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
defparam \Selector5~0 .lut_mask = 16'h88F8;
defparam \Selector5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_state~0 (
	.dataa(out_rsp_data_0),
	.datab(\current_state.STATE_POLL_RSP~q ),
	.datac(\busy~0_combout ),
	.datad(\current_state.STATE_STATUS_RSP~q ),
	.cin(gnd),
	.combout(\next_state~0_combout ),
	.cout());
defparam \next_state~0 .lut_mask = 16'hAAC0;
defparam \next_state~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~0 (
	.dataa(\always0~0_combout ),
	.datab(\current_state.STATE_STATUS_RSP~q ),
	.datac(\next_state~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'h8080;
defparam \Selector1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \fifo_in_valid~0 (
	.dataa(\mem_wr_combi~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avst_fifo_inst|avst_fifo|full~q ),
	.cin(gnd),
	.combout(\fifo_in_valid~0_combout ),
	.cout());
defparam \fifo_in_valid~0 .lut_mask = 16'h00AA;
defparam \fifo_in_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector10~0 (
	.dataa(hold_waitrequest1),
	.datab(avl_mem_read),
	.datac(gnd),
	.datad(\current_state.STATE_IDLE~q ),
	.cin(gnd),
	.combout(\Selector10~0_combout ),
	.cout());
defparam \Selector10~0 .lut_mask = 16'h0088;
defparam \Selector10~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~1 (
	.dataa(\Equal2~1_combout ),
	.datab(\fifo_in_valid~0_combout ),
	.datac(\current_state.STATE_IDLE~q ),
	.datad(\Selector10~0_combout ),
	.cin(gnd),
	.combout(\Selector1~1_combout ),
	.cout());
defparam \Selector1~1 .lut_mask = 16'h0008;
defparam \Selector1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~2 (
	.dataa(\Selector1~0_combout ),
	.datab(\Selector1~1_combout ),
	.datac(current_stateSTATE_STATUS_CMD),
	.datad(sink0_ready),
	.cin(gnd),
	.combout(\Selector1~2_combout ),
	.cout());
defparam \Selector1~2 .lut_mask = 16'hEEFE;
defparam \Selector1~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector7~0 (
	.dataa(\always0~0_combout ),
	.datab(current_stateSTATE_WR_DATA),
	.datac(\current_state.STATE_POLL_RSP~q ),
	.datad(\next_state~0_combout ),
	.cin(gnd),
	.combout(\Selector7~0_combout ),
	.cout());
defparam \Selector7~0 .lut_mask = 16'hA888;
defparam \Selector7~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector7~1 (
	.dataa(\Selector7~0_combout ),
	.datab(current_stateSTATE_POLL_CMD),
	.datac(gnd),
	.datad(sink0_ready),
	.cin(gnd),
	.combout(\Selector7~1_combout ),
	.cout());
defparam \Selector7~1 .lut_mask = 16'hAAEE;
defparam \Selector7~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector10~1 (
	.dataa(\Selector10~0_combout ),
	.datab(current_stateSTATE_READ_CMD),
	.datac(\current_state.STATE_IDLE~q ),
	.datad(sink0_ready),
	.cin(gnd),
	.combout(\Selector10~1_combout ),
	.cout());
defparam \Selector10~1 .lut_mask = 16'h0ACE;
defparam \Selector10~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector6~0 (
	.dataa(current_stateSTATE_WR_CMD),
	.datab(sink0_ready),
	.datac(current_stateSTATE_WR_DATA),
	.datad(\always0~0_combout ),
	.cin(gnd),
	.combout(\Selector6~0_combout ),
	.cout());
defparam \Selector6~0 .lut_mask = 16'h88F8;
defparam \Selector6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always10~2 (
	.dataa(\mem_wr_combi~0_combout ),
	.datab(\avst_fifo_inst|avst_fifo|full~q ),
	.datac(\Selector10~0_combout ),
	.datad(\Equal2~1_combout ),
	.cin(gnd),
	.combout(\always10~2_combout ),
	.cout());
defparam \always10~2 .lut_mask = 16'hF2F0;
defparam \always10~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_byteenable_reg[0]~0 (
	.dataa(mem_burstcount[2]),
	.datab(mem_burstcount[1]),
	.datac(mem_burstcount[4]),
	.datad(mem_burstcount[3]),
	.cin(gnd),
	.combout(\mem_byteenable_reg[0]~0_combout ),
	.cout());
defparam \mem_byteenable_reg[0]~0 .lut_mask = 16'h0001;
defparam \mem_byteenable_reg[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_byteenable_reg[0]~1 (
	.dataa(\mem_byteenable_reg[0]~0_combout ),
	.datab(gnd),
	.datac(mem_burstcount[6]),
	.datad(mem_burstcount[5]),
	.cin(gnd),
	.combout(\mem_byteenable_reg[0]~1_combout ),
	.cout());
defparam \mem_byteenable_reg[0]~1 .lut_mask = 16'h000A;
defparam \mem_byteenable_reg[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \is_burst_reg~0 (
	.dataa(is_burst_reg1),
	.datab(gnd),
	.datac(\always10~2_combout ),
	.datad(\mem_byteenable_reg[0]~1_combout ),
	.cin(gnd),
	.combout(\is_burst_reg~0_combout ),
	.cout());
defparam \is_burst_reg~0 .lut_mask = 16'h0AFA;
defparam \is_burst_reg~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_byteenable_reg~2 (
	.dataa(avl_mem_byteenable_0),
	.datab(mem_burstcount[0]),
	.datac(\mem_wr_combi~0_combout ),
	.datad(\mem_byteenable_reg[0]~1_combout ),
	.cin(gnd),
	.combout(\mem_byteenable_reg~2_combout ),
	.cout());
defparam \mem_byteenable_reg~2 .lut_mask = 16'hBFFF;
defparam \mem_byteenable_reg~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_byteenable_reg[0]~3 (
	.dataa(\Equal0~0_combout ),
	.datab(avl_mem_write),
	.datac(avl_mem_read),
	.datad(mem_waitrequest),
	.cin(gnd),
	.combout(\mem_byteenable_reg[0]~3_combout ),
	.cout());
defparam \mem_byteenable_reg[0]~3 .lut_mask = 16'hF400;
defparam \mem_byteenable_reg[0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_byteenable_reg~4 (
	.dataa(avl_mem_byteenable_3),
	.datab(mem_burstcount[0]),
	.datac(\mem_wr_combi~0_combout ),
	.datad(\mem_byteenable_reg[0]~1_combout ),
	.cin(gnd),
	.combout(\mem_byteenable_reg~4_combout ),
	.cout());
defparam \mem_byteenable_reg~4 .lut_mask = 16'hBFFF;
defparam \mem_byteenable_reg~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_byteenable_reg~5 (
	.dataa(avl_mem_byteenable_2),
	.datab(mem_burstcount[0]),
	.datac(\mem_wr_combi~0_combout ),
	.datad(\mem_byteenable_reg[0]~1_combout ),
	.cin(gnd),
	.combout(\mem_byteenable_reg~5_combout ),
	.cout());
defparam \mem_byteenable_reg~5 .lut_mask = 16'hBFFF;
defparam \mem_byteenable_reg~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_byteenable_reg~6 (
	.dataa(avl_mem_byteenable_1),
	.datab(mem_burstcount[0]),
	.datac(\mem_wr_combi~0_combout ),
	.datad(\mem_byteenable_reg[0]~1_combout ),
	.cin(gnd),
	.combout(\mem_byteenable_reg~6_combout ),
	.cout());
defparam \mem_byteenable_reg~6 .lut_mask = 16'hBFFF;
defparam \mem_byteenable_reg~6 .sum_lutc_input = "datac";

dffeas \mem_write_data_reg[11] (
	.clk(clk_clk),
	.d(avl_mem_writedata_11),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(\mem_write_data_reg[11]~q ),
	.prn(vcc));
defparam \mem_write_data_reg[11] .is_wysiwyg = "true";
defparam \mem_write_data_reg[11] .power_up = "low";

cycloneive_lcell_comb \cmd_data[11]~4 (
	.dataa(mem_byteenable_reg_3),
	.datab(mem_byteenable_reg_2),
	.datac(mem_write_data_reg_27),
	.datad(mem_byteenable_reg_0),
	.cin(gnd),
	.combout(\cmd_data[11]~4_combout ),
	.cout());
defparam \cmd_data[11]~4 .lut_mask = 16'h0080;
defparam \cmd_data[11]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(mem_byteenable_reg_3),
	.datad(mem_byteenable_reg_2),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout());
defparam \Add1~0 .lut_mask = 16'h0FF0;
defparam \Add1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[8]~5 (
	.dataa(mem_byteenable_reg_1),
	.datab(is_burst_reg1),
	.datac(\Add1~0_combout ),
	.datad(current_stateSTATE_WR_DATA),
	.cin(gnd),
	.combout(\cmd_data[8]~5_combout ),
	.cout());
defparam \cmd_data[8]~5 .lut_mask = 16'h02FF;
defparam \cmd_data[8]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[8]~88 (
	.dataa(is_burst_reg1),
	.datab(current_stateSTATE_WR_DATA),
	.datac(mem_byteenable_reg_0),
	.datad(\cmd_data[8]~5_combout ),
	.cin(gnd),
	.combout(\cmd_data[8]~88_combout ),
	.cout());
defparam \cmd_data[8]~88 .lut_mask = 16'h4044;
defparam \cmd_data[8]~88 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector17~0 (
	.dataa(gnd),
	.datab(current_stateSTATE_WR_CMD),
	.datac(\current_state.STATE_WRENABLE_CMD~q ),
	.datad(WideOr13),
	.cin(gnd),
	.combout(\Selector17~0_combout ),
	.cout());
defparam \Selector17~0 .lut_mask = 16'h0003;
defparam \Selector17~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[8]~6 (
	.dataa(is_burst_reg1),
	.datab(gnd),
	.datac(gnd),
	.datad(current_stateSTATE_WR_DATA),
	.cin(gnd),
	.combout(\cmd_data[8]~6_combout ),
	.cout());
defparam \cmd_data[8]~6 .lut_mask = 16'hAAFF;
defparam \cmd_data[8]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[11]~7 (
	.dataa(\Selector17~0_combout ),
	.datab(\avst_fifo_inst|avst_fifo|out_payload[11]~q ),
	.datac(\cmd_data[8]~6_combout ),
	.datad(\cmd_data[8]~5_combout ),
	.cin(gnd),
	.combout(\cmd_data[11]~7_combout ),
	.cout());
defparam \cmd_data[11]~7 .lut_mask = 16'hA0CF;
defparam \cmd_data[11]~7 .sum_lutc_input = "datac";

dffeas \mem_write_data_reg[10] (
	.clk(clk_clk),
	.d(avl_mem_writedata_10),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(\mem_write_data_reg[10]~q ),
	.prn(vcc));
defparam \mem_write_data_reg[10] .is_wysiwyg = "true";
defparam \mem_write_data_reg[10] .power_up = "low";

cycloneive_lcell_comb \cmd_data[10]~8 (
	.dataa(mem_byteenable_reg_3),
	.datab(mem_byteenable_reg_2),
	.datac(mem_write_data_reg_26),
	.datad(mem_byteenable_reg_0),
	.cin(gnd),
	.combout(\cmd_data[10]~8_combout ),
	.cout());
defparam \cmd_data[10]~8 .lut_mask = 16'h0080;
defparam \cmd_data[10]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[10]~9 (
	.dataa(current_stateSTATE_WR_CMD),
	.datab(\avst_fifo_inst|avst_fifo|out_payload[10]~q ),
	.datac(\cmd_data[8]~6_combout ),
	.datad(\cmd_data[8]~5_combout ),
	.cin(gnd),
	.combout(\cmd_data[10]~9_combout ),
	.cout());
defparam \cmd_data[10]~9 .lut_mask = 16'hA0CF;
defparam \cmd_data[10]~9 .sum_lutc_input = "datac";

dffeas \mem_write_data_reg[8] (
	.clk(clk_clk),
	.d(avl_mem_writedata_8),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(\mem_write_data_reg[8]~q ),
	.prn(vcc));
defparam \mem_write_data_reg[8] .is_wysiwyg = "true";
defparam \mem_write_data_reg[8] .power_up = "low";

cycloneive_lcell_comb \cmd_data[8]~10 (
	.dataa(mem_byteenable_reg_3),
	.datab(mem_byteenable_reg_2),
	.datac(mem_write_data_reg_24),
	.datad(mem_byteenable_reg_0),
	.cin(gnd),
	.combout(\cmd_data[8]~10_combout ),
	.cout());
defparam \cmd_data[8]~10 .lut_mask = 16'h0080;
defparam \cmd_data[8]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[8]~11 (
	.dataa(Selector20),
	.datab(\avst_fifo_inst|avst_fifo|out_payload[8]~q ),
	.datac(\cmd_data[8]~6_combout ),
	.datad(\cmd_data[8]~5_combout ),
	.cin(gnd),
	.combout(\cmd_data[8]~11_combout ),
	.cout());
defparam \cmd_data[8]~11 .lut_mask = 16'h50CF;
defparam \cmd_data[8]~11 .sum_lutc_input = "datac";

dffeas \mem_write_data_reg[13] (
	.clk(clk_clk),
	.d(avl_mem_writedata_13),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(\mem_write_data_reg[13]~q ),
	.prn(vcc));
defparam \mem_write_data_reg[13] .is_wysiwyg = "true";
defparam \mem_write_data_reg[13] .power_up = "low";

cycloneive_lcell_comb \cmd_data[13]~12 (
	.dataa(mem_byteenable_reg_3),
	.datab(mem_byteenable_reg_2),
	.datac(mem_write_data_reg_29),
	.datad(mem_byteenable_reg_0),
	.cin(gnd),
	.combout(\cmd_data[13]~12_combout ),
	.cout());
defparam \cmd_data[13]~12 .lut_mask = 16'h0080;
defparam \cmd_data[13]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector15~0 (
	.dataa(current_stateSTATE_WR_CMD),
	.datab(csr_rd_inst_data_8),
	.datac(current_stateSTATE_READ_CMD),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector15~0_combout ),
	.cout());
defparam \Selector15~0 .lut_mask = 16'hEAEA;
defparam \Selector15~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[13]~13 (
	.dataa(\Selector15~0_combout ),
	.datab(\avst_fifo_inst|avst_fifo|out_payload[13]~q ),
	.datac(\cmd_data[8]~6_combout ),
	.datad(\cmd_data[8]~5_combout ),
	.cin(gnd),
	.combout(\cmd_data[13]~13_combout ),
	.cout());
defparam \cmd_data[13]~13 .lut_mask = 16'hA0CF;
defparam \cmd_data[13]~13 .sum_lutc_input = "datac";

dffeas \mem_write_data_reg[15] (
	.clk(clk_clk),
	.d(avl_mem_writedata_15),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(\mem_write_data_reg[15]~q ),
	.prn(vcc));
defparam \mem_write_data_reg[15] .is_wysiwyg = "true";
defparam \mem_write_data_reg[15] .power_up = "low";

cycloneive_lcell_comb \cmd_data[15]~14 (
	.dataa(mem_byteenable_reg_3),
	.datab(mem_byteenable_reg_2),
	.datac(mem_write_data_reg_31),
	.datad(mem_byteenable_reg_0),
	.cin(gnd),
	.combout(\cmd_data[15]~14_combout ),
	.cout());
defparam \cmd_data[15]~14 .lut_mask = 16'h0080;
defparam \cmd_data[15]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[14]~15 (
	.dataa(current_stateSTATE_WR_DATA),
	.datab(is_burst_reg1),
	.datac(mem_byteenable_reg_1),
	.datad(\Add1~0_combout ),
	.cin(gnd),
	.combout(\cmd_data[14]~15_combout ),
	.cout());
defparam \cmd_data[14]~15 .lut_mask = 16'h88A8;
defparam \cmd_data[14]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[14]~89 (
	.dataa(is_burst_reg1),
	.datab(current_stateSTATE_WR_DATA),
	.datac(mem_byteenable_reg_0),
	.datad(\cmd_data[14]~15_combout ),
	.cin(gnd),
	.combout(\cmd_data[14]~89_combout ),
	.cout());
defparam \cmd_data[14]~89 .lut_mask = 16'h4044;
defparam \cmd_data[14]~89 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[15]~16 (
	.dataa(csr_rd_inst_data_10),
	.datab(current_stateSTATE_READ_CMD),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\cmd_data[15]~16_combout ),
	.cout());
defparam \cmd_data[15]~16 .lut_mask = 16'h8888;
defparam \cmd_data[15]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[15]~17 (
	.dataa(\avst_fifo_inst|avst_fifo|out_payload[15]~q ),
	.datab(\cmd_data[15]~16_combout ),
	.datac(\cmd_data[8]~6_combout ),
	.datad(\cmd_data[14]~15_combout ),
	.cin(gnd),
	.combout(\cmd_data[15]~17_combout ),
	.cout());
defparam \cmd_data[15]~17 .lut_mask = 16'hA0CF;
defparam \cmd_data[15]~17 .sum_lutc_input = "datac";

dffeas \mem_write_data_reg[14] (
	.clk(clk_clk),
	.d(avl_mem_writedata_14),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(\mem_write_data_reg[14]~q ),
	.prn(vcc));
defparam \mem_write_data_reg[14] .is_wysiwyg = "true";
defparam \mem_write_data_reg[14] .power_up = "low";

cycloneive_lcell_comb \cmd_data[14]~18 (
	.dataa(mem_write_data_reg_30),
	.datab(mem_byteenable_reg_3),
	.datac(mem_byteenable_reg_2),
	.datad(mem_byteenable_reg_0),
	.cin(gnd),
	.combout(\cmd_data[14]~18_combout ),
	.cout());
defparam \cmd_data[14]~18 .lut_mask = 16'h0080;
defparam \cmd_data[14]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[14]~19 (
	.dataa(csr_rd_inst_data_9),
	.datab(current_stateSTATE_READ_CMD),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\cmd_data[14]~19_combout ),
	.cout());
defparam \cmd_data[14]~19 .lut_mask = 16'h8888;
defparam \cmd_data[14]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[14]~20 (
	.dataa(\avst_fifo_inst|avst_fifo|out_payload[14]~q ),
	.datab(\cmd_data[14]~19_combout ),
	.datac(\cmd_data[8]~6_combout ),
	.datad(\cmd_data[14]~15_combout ),
	.cin(gnd),
	.combout(\cmd_data[14]~20_combout ),
	.cout());
defparam \cmd_data[14]~20 .lut_mask = 16'hA0CF;
defparam \cmd_data[14]~20 .sum_lutc_input = "datac";

dffeas \mem_write_data_reg[9] (
	.clk(clk_clk),
	.d(avl_mem_writedata_9),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(\mem_write_data_reg[9]~q ),
	.prn(vcc));
defparam \mem_write_data_reg[9] .is_wysiwyg = "true";
defparam \mem_write_data_reg[9] .power_up = "low";

cycloneive_lcell_comb \cmd_data[9]~21 (
	.dataa(mem_byteenable_reg_3),
	.datab(mem_byteenable_reg_2),
	.datac(mem_write_data_reg_25),
	.datad(mem_byteenable_reg_0),
	.cin(gnd),
	.combout(\cmd_data[9]~21_combout ),
	.cout());
defparam \cmd_data[9]~21 .lut_mask = 16'h0080;
defparam \cmd_data[9]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector19~0 (
	.dataa(csr_control_data_8),
	.datab(current_stateSTATE_WR_CMD),
	.datac(current_stateSTATE_READ_CMD),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector19~0_combout ),
	.cout());
defparam \Selector19~0 .lut_mask = 16'hA8A8;
defparam \Selector19~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[9]~22 (
	.dataa(\Selector19~0_combout ),
	.datab(\avst_fifo_inst|avst_fifo|out_payload[9]~q ),
	.datac(\cmd_data[8]~6_combout ),
	.datad(\cmd_data[8]~5_combout ),
	.cin(gnd),
	.combout(\cmd_data[9]~22_combout ),
	.cout());
defparam \cmd_data[9]~22 .lut_mask = 16'hA0CF;
defparam \cmd_data[9]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[0]~23 (
	.dataa(csr_wr_inst_data_0),
	.datab(current_stateSTATE_STATUS_CMD),
	.datac(gnd),
	.datad(current_stateSTATE_WR_CMD),
	.cin(gnd),
	.combout(\cmd_data[0]~23_combout ),
	.cout());
defparam \cmd_data[0]~23 .lut_mask = 16'hAACC;
defparam \cmd_data[0]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[2]~24 (
	.dataa(current_stateSTATE_WR_DATA),
	.datab(current_stateSTATE_READ_CMD),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\cmd_data[2]~24_combout ),
	.cout());
defparam \cmd_data[2]~24 .lut_mask = 16'hEEEE;
defparam \cmd_data[2]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[2]~25 (
	.dataa(mem_byteenable_reg_3),
	.datab(mem_byteenable_reg_2),
	.datac(mem_byteenable_reg_0),
	.datad(mem_byteenable_reg_1),
	.cin(gnd),
	.combout(\cmd_data[2]~25_combout ),
	.cout());
defparam \cmd_data[2]~25 .lut_mask = 16'h2AEE;
defparam \cmd_data[2]~25 .sum_lutc_input = "datac";

dffeas \mem_write_data_reg[0] (
	.clk(clk_clk),
	.d(avl_mem_writedata_0),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(\mem_write_data_reg[0]~q ),
	.prn(vcc));
defparam \mem_write_data_reg[0] .is_wysiwyg = "true";
defparam \mem_write_data_reg[0] .power_up = "low";

cycloneive_lcell_comb \cmd_data[2]~26 (
	.dataa(mem_byteenable_reg_1),
	.datab(mem_byteenable_reg_3),
	.datac(mem_byteenable_reg_0),
	.datad(mem_byteenable_reg_2),
	.cin(gnd),
	.combout(\cmd_data[2]~26_combout ),
	.cout());
defparam \cmd_data[2]~26 .lut_mask = 16'h2ACF;
defparam \cmd_data[2]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[0]~27 (
	.dataa(mem_write_data_reg_16),
	.datab(\mem_write_data_reg[0]~q ),
	.datac(\cmd_data[2]~26_combout ),
	.datad(\cmd_data[2]~25_combout ),
	.cin(gnd),
	.combout(\cmd_data[0]~27_combout ),
	.cout());
defparam \cmd_data[0]~27 .lut_mask = 16'h0AFC;
defparam \cmd_data[0]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[2]~28 (
	.dataa(mem_byteenable_reg_0),
	.datab(mem_byteenable_reg_1),
	.datac(mem_byteenable_reg_2),
	.datad(mem_byteenable_reg_3),
	.cin(gnd),
	.combout(\cmd_data[2]~28_combout ),
	.cout());
defparam \cmd_data[2]~28 .lut_mask = 16'h03C5;
defparam \cmd_data[2]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[0]~29 (
	.dataa(gnd),
	.datab(\mem_write_data_reg[8]~q ),
	.datac(mem_byteenable_reg_2),
	.datad(gnd),
	.cin(gnd),
	.combout(\cmd_data[0]~29_combout ),
	.cout());
defparam \cmd_data[0]~29 .lut_mask = 16'h0C0C;
defparam \cmd_data[0]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[0]~30 (
	.dataa(mem_write_data_reg_24),
	.datab(\cmd_data[2]~28_combout ),
	.datac(\cmd_data[0]~29_combout ),
	.datad(\cmd_data[0]~27_combout ),
	.cin(gnd),
	.combout(\cmd_data[0]~30_combout ),
	.cout());
defparam \cmd_data[0]~30 .lut_mask = 16'h0C88;
defparam \cmd_data[0]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[0]~31 (
	.dataa(mem_byteenable_reg_0),
	.datab(\cmd_data[2]~25_combout ),
	.datac(\cmd_data[0]~27_combout ),
	.datad(\cmd_data[0]~30_combout ),
	.cin(gnd),
	.combout(\cmd_data[0]~31_combout ),
	.cout());
defparam \cmd_data[0]~31 .lut_mask = 16'h0570;
defparam \cmd_data[0]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[2]~32 (
	.dataa(mem_byteenable_reg_0),
	.datab(mem_byteenable_reg_3),
	.datac(mem_byteenable_reg_2),
	.datad(mem_byteenable_reg_1),
	.cin(gnd),
	.combout(\cmd_data[2]~32_combout ),
	.cout());
defparam \cmd_data[2]~32 .lut_mask = 16'hBFFE;
defparam \cmd_data[2]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[2]~33 (
	.dataa(\cmd_data[2]~32_combout ),
	.datab(current_stateSTATE_READ_CMD),
	.datac(gnd),
	.datad(current_stateSTATE_WR_DATA),
	.cin(gnd),
	.combout(\cmd_data[2]~33_combout ),
	.cout());
defparam \cmd_data[2]~33 .lut_mask = 16'hAACC;
defparam \cmd_data[2]~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[2]~34 (
	.dataa(current_stateSTATE_POLL_CMD),
	.datab(current_stateSTATE_READ_CMD),
	.datac(gnd),
	.datad(current_stateSTATE_WR_DATA),
	.cin(gnd),
	.combout(\cmd_data[2]~34_combout ),
	.cout());
defparam \cmd_data[2]~34 .lut_mask = 16'h00EE;
defparam \cmd_data[2]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[0]~35 (
	.dataa(\cmd_data[0]~31_combout ),
	.datab(csr_rd_inst_data_0),
	.datac(\cmd_data[2]~33_combout ),
	.datad(\cmd_data[2]~34_combout ),
	.cin(gnd),
	.combout(\cmd_data[0]~35_combout ),
	.cout());
defparam \cmd_data[0]~35 .lut_mask = 16'h3FA0;
defparam \cmd_data[0]~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[4]~37 (
	.dataa(csr_wr_inst_data_4),
	.datab(current_stateSTATE_WR_CMD),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\cmd_data[4]~37_combout ),
	.cout());
defparam \cmd_data[4]~37 .lut_mask = 16'h8888;
defparam \cmd_data[4]~37 .sum_lutc_input = "datac";

dffeas \mem_write_data_reg[4] (
	.clk(clk_clk),
	.d(avl_mem_writedata_4),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(\mem_write_data_reg[4]~q ),
	.prn(vcc));
defparam \mem_write_data_reg[4] .is_wysiwyg = "true";
defparam \mem_write_data_reg[4] .power_up = "low";

cycloneive_lcell_comb \cmd_data[4]~38 (
	.dataa(mem_write_data_reg_20),
	.datab(\mem_write_data_reg[4]~q ),
	.datac(\cmd_data[2]~26_combout ),
	.datad(\cmd_data[2]~25_combout ),
	.cin(gnd),
	.combout(\cmd_data[4]~38_combout ),
	.cout());
defparam \cmd_data[4]~38 .lut_mask = 16'h0AFC;
defparam \cmd_data[4]~38 .sum_lutc_input = "datac";

dffeas \mem_write_data_reg[12] (
	.clk(clk_clk),
	.d(avl_mem_writedata_12),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(\mem_write_data_reg[12]~q ),
	.prn(vcc));
defparam \mem_write_data_reg[12] .is_wysiwyg = "true";
defparam \mem_write_data_reg[12] .power_up = "low";

cycloneive_lcell_comb \cmd_data[4]~39 (
	.dataa(gnd),
	.datab(\mem_write_data_reg[12]~q ),
	.datac(mem_byteenable_reg_2),
	.datad(gnd),
	.cin(gnd),
	.combout(\cmd_data[4]~39_combout ),
	.cout());
defparam \cmd_data[4]~39 .lut_mask = 16'h0C0C;
defparam \cmd_data[4]~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[4]~40 (
	.dataa(mem_write_data_reg_28),
	.datab(\cmd_data[2]~28_combout ),
	.datac(\cmd_data[4]~39_combout ),
	.datad(\cmd_data[4]~38_combout ),
	.cin(gnd),
	.combout(\cmd_data[4]~40_combout ),
	.cout());
defparam \cmd_data[4]~40 .lut_mask = 16'h0C88;
defparam \cmd_data[4]~40 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[4]~41 (
	.dataa(mem_byteenable_reg_0),
	.datab(\cmd_data[2]~25_combout ),
	.datac(\cmd_data[4]~38_combout ),
	.datad(\cmd_data[4]~40_combout ),
	.cin(gnd),
	.combout(\cmd_data[4]~41_combout ),
	.cout());
defparam \cmd_data[4]~41 .lut_mask = 16'h0570;
defparam \cmd_data[4]~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[4]~42 (
	.dataa(\cmd_data[4]~41_combout ),
	.datab(csr_rd_inst_data_4),
	.datac(\cmd_data[2]~33_combout ),
	.datad(\cmd_data[2]~34_combout ),
	.cin(gnd),
	.combout(\cmd_data[4]~42_combout ),
	.cout());
defparam \cmd_data[4]~42 .lut_mask = 16'hCFA0;
defparam \cmd_data[4]~42 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[2]~44 (
	.dataa(csr_wr_inst_data_2),
	.datab(current_stateSTATE_STATUS_CMD),
	.datac(\current_state.STATE_WRENABLE_CMD~q ),
	.datad(current_stateSTATE_WR_CMD),
	.cin(gnd),
	.combout(\cmd_data[2]~44_combout ),
	.cout());
defparam \cmd_data[2]~44 .lut_mask = 16'hAAFC;
defparam \cmd_data[2]~44 .sum_lutc_input = "datac";

dffeas \mem_write_data_reg[2] (
	.clk(clk_clk),
	.d(avl_mem_writedata_2),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(\mem_write_data_reg[2]~q ),
	.prn(vcc));
defparam \mem_write_data_reg[2] .is_wysiwyg = "true";
defparam \mem_write_data_reg[2] .power_up = "low";

cycloneive_lcell_comb \cmd_data[2]~45 (
	.dataa(mem_write_data_reg_18),
	.datab(\mem_write_data_reg[2]~q ),
	.datac(\cmd_data[2]~26_combout ),
	.datad(\cmd_data[2]~25_combout ),
	.cin(gnd),
	.combout(\cmd_data[2]~45_combout ),
	.cout());
defparam \cmd_data[2]~45 .lut_mask = 16'h0AFC;
defparam \cmd_data[2]~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[2]~46 (
	.dataa(gnd),
	.datab(\mem_write_data_reg[10]~q ),
	.datac(mem_byteenable_reg_2),
	.datad(gnd),
	.cin(gnd),
	.combout(\cmd_data[2]~46_combout ),
	.cout());
defparam \cmd_data[2]~46 .lut_mask = 16'h0C0C;
defparam \cmd_data[2]~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[2]~47 (
	.dataa(mem_write_data_reg_26),
	.datab(\cmd_data[2]~28_combout ),
	.datac(\cmd_data[2]~46_combout ),
	.datad(\cmd_data[2]~45_combout ),
	.cin(gnd),
	.combout(\cmd_data[2]~47_combout ),
	.cout());
defparam \cmd_data[2]~47 .lut_mask = 16'h0C88;
defparam \cmd_data[2]~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[2]~48 (
	.dataa(mem_byteenable_reg_0),
	.datab(\cmd_data[2]~25_combout ),
	.datac(\cmd_data[2]~45_combout ),
	.datad(\cmd_data[2]~47_combout ),
	.cin(gnd),
	.combout(\cmd_data[2]~48_combout ),
	.cout());
defparam \cmd_data[2]~48 .lut_mask = 16'h0570;
defparam \cmd_data[2]~48 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[2]~49 (
	.dataa(\cmd_data[2]~48_combout ),
	.datab(csr_rd_inst_data_2),
	.datac(\cmd_data[2]~33_combout ),
	.datad(\cmd_data[2]~34_combout ),
	.cin(gnd),
	.combout(\cmd_data[2]~49_combout ),
	.cout());
defparam \cmd_data[2]~49 .lut_mask = 16'hCFA0;
defparam \cmd_data[2]~49 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[1]~51 (
	.dataa(\current_state.STATE_WRENABLE_CMD~q ),
	.datab(gnd),
	.datac(current_stateSTATE_WR_CMD),
	.datad(csr_wr_inst_data_1),
	.cin(gnd),
	.combout(\cmd_data[1]~51_combout ),
	.cout());
defparam \cmd_data[1]~51 .lut_mask = 16'h0AFA;
defparam \cmd_data[1]~51 .sum_lutc_input = "datac";

dffeas \mem_write_data_reg[1] (
	.clk(clk_clk),
	.d(avl_mem_writedata_1),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(\mem_write_data_reg[1]~q ),
	.prn(vcc));
defparam \mem_write_data_reg[1] .is_wysiwyg = "true";
defparam \mem_write_data_reg[1] .power_up = "low";

cycloneive_lcell_comb \cmd_data[1]~52 (
	.dataa(mem_write_data_reg_17),
	.datab(\mem_write_data_reg[1]~q ),
	.datac(\cmd_data[2]~26_combout ),
	.datad(\cmd_data[2]~25_combout ),
	.cin(gnd),
	.combout(\cmd_data[1]~52_combout ),
	.cout());
defparam \cmd_data[1]~52 .lut_mask = 16'h0AFC;
defparam \cmd_data[1]~52 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[1]~53 (
	.dataa(gnd),
	.datab(\mem_write_data_reg[9]~q ),
	.datac(mem_byteenable_reg_2),
	.datad(gnd),
	.cin(gnd),
	.combout(\cmd_data[1]~53_combout ),
	.cout());
defparam \cmd_data[1]~53 .lut_mask = 16'h0C0C;
defparam \cmd_data[1]~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[1]~54 (
	.dataa(mem_write_data_reg_25),
	.datab(\cmd_data[2]~28_combout ),
	.datac(\cmd_data[1]~53_combout ),
	.datad(\cmd_data[1]~52_combout ),
	.cin(gnd),
	.combout(\cmd_data[1]~54_combout ),
	.cout());
defparam \cmd_data[1]~54 .lut_mask = 16'h0C88;
defparam \cmd_data[1]~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[1]~55 (
	.dataa(mem_byteenable_reg_0),
	.datab(\cmd_data[2]~25_combout ),
	.datac(\cmd_data[1]~52_combout ),
	.datad(\cmd_data[1]~54_combout ),
	.cin(gnd),
	.combout(\cmd_data[1]~55_combout ),
	.cout());
defparam \cmd_data[1]~55 .lut_mask = 16'h0570;
defparam \cmd_data[1]~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[1]~56 (
	.dataa(\cmd_data[1]~55_combout ),
	.datab(csr_rd_inst_data_1),
	.datac(\cmd_data[2]~33_combout ),
	.datad(\cmd_data[2]~34_combout ),
	.cin(gnd),
	.combout(\cmd_data[1]~56_combout ),
	.cout());
defparam \cmd_data[1]~56 .lut_mask = 16'h3FA0;
defparam \cmd_data[1]~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[3]~58 (
	.dataa(csr_wr_inst_data_3),
	.datab(current_stateSTATE_WR_CMD),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\cmd_data[3]~58_combout ),
	.cout());
defparam \cmd_data[3]~58 .lut_mask = 16'h8888;
defparam \cmd_data[3]~58 .sum_lutc_input = "datac";

dffeas \mem_write_data_reg[3] (
	.clk(clk_clk),
	.d(avl_mem_writedata_3),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(\mem_write_data_reg[3]~q ),
	.prn(vcc));
defparam \mem_write_data_reg[3] .is_wysiwyg = "true";
defparam \mem_write_data_reg[3] .power_up = "low";

cycloneive_lcell_comb \cmd_data[3]~59 (
	.dataa(mem_write_data_reg_19),
	.datab(\mem_write_data_reg[3]~q ),
	.datac(\cmd_data[2]~26_combout ),
	.datad(\cmd_data[2]~25_combout ),
	.cin(gnd),
	.combout(\cmd_data[3]~59_combout ),
	.cout());
defparam \cmd_data[3]~59 .lut_mask = 16'h0AFC;
defparam \cmd_data[3]~59 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[3]~60 (
	.dataa(gnd),
	.datab(\mem_write_data_reg[11]~q ),
	.datac(mem_byteenable_reg_2),
	.datad(gnd),
	.cin(gnd),
	.combout(\cmd_data[3]~60_combout ),
	.cout());
defparam \cmd_data[3]~60 .lut_mask = 16'h0C0C;
defparam \cmd_data[3]~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[3]~61 (
	.dataa(mem_write_data_reg_27),
	.datab(\cmd_data[2]~28_combout ),
	.datac(\cmd_data[3]~60_combout ),
	.datad(\cmd_data[3]~59_combout ),
	.cin(gnd),
	.combout(\cmd_data[3]~61_combout ),
	.cout());
defparam \cmd_data[3]~61 .lut_mask = 16'h0C88;
defparam \cmd_data[3]~61 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[3]~62 (
	.dataa(mem_byteenable_reg_0),
	.datab(\cmd_data[2]~25_combout ),
	.datac(\cmd_data[3]~59_combout ),
	.datad(\cmd_data[3]~61_combout ),
	.cin(gnd),
	.combout(\cmd_data[3]~62_combout ),
	.cout());
defparam \cmd_data[3]~62 .lut_mask = 16'h0570;
defparam \cmd_data[3]~62 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[3]~63 (
	.dataa(\cmd_data[3]~62_combout ),
	.datab(csr_rd_inst_data_3),
	.datac(\cmd_data[2]~33_combout ),
	.datad(\cmd_data[2]~34_combout ),
	.cin(gnd),
	.combout(\cmd_data[3]~63_combout ),
	.cout());
defparam \cmd_data[3]~63 .lut_mask = 16'hCFA0;
defparam \cmd_data[3]~63 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[5]~65 (
	.dataa(csr_wr_inst_data_5),
	.datab(current_stateSTATE_WR_CMD),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\cmd_data[5]~65_combout ),
	.cout());
defparam \cmd_data[5]~65 .lut_mask = 16'h8888;
defparam \cmd_data[5]~65 .sum_lutc_input = "datac";

dffeas \mem_write_data_reg[5] (
	.clk(clk_clk),
	.d(avl_mem_writedata_5),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(\mem_write_data_reg[5]~q ),
	.prn(vcc));
defparam \mem_write_data_reg[5] .is_wysiwyg = "true";
defparam \mem_write_data_reg[5] .power_up = "low";

cycloneive_lcell_comb \cmd_data[5]~66 (
	.dataa(mem_write_data_reg_21),
	.datab(\mem_write_data_reg[5]~q ),
	.datac(\cmd_data[2]~26_combout ),
	.datad(\cmd_data[2]~25_combout ),
	.cin(gnd),
	.combout(\cmd_data[5]~66_combout ),
	.cout());
defparam \cmd_data[5]~66 .lut_mask = 16'h0AFC;
defparam \cmd_data[5]~66 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[5]~67 (
	.dataa(gnd),
	.datab(\mem_write_data_reg[13]~q ),
	.datac(mem_byteenable_reg_2),
	.datad(gnd),
	.cin(gnd),
	.combout(\cmd_data[5]~67_combout ),
	.cout());
defparam \cmd_data[5]~67 .lut_mask = 16'h0C0C;
defparam \cmd_data[5]~67 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[5]~68 (
	.dataa(mem_write_data_reg_29),
	.datab(\cmd_data[2]~28_combout ),
	.datac(\cmd_data[5]~67_combout ),
	.datad(\cmd_data[5]~66_combout ),
	.cin(gnd),
	.combout(\cmd_data[5]~68_combout ),
	.cout());
defparam \cmd_data[5]~68 .lut_mask = 16'h0C88;
defparam \cmd_data[5]~68 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[5]~69 (
	.dataa(mem_byteenable_reg_0),
	.datab(\cmd_data[2]~25_combout ),
	.datac(\cmd_data[5]~66_combout ),
	.datad(\cmd_data[5]~68_combout ),
	.cin(gnd),
	.combout(\cmd_data[5]~69_combout ),
	.cout());
defparam \cmd_data[5]~69 .lut_mask = 16'h0570;
defparam \cmd_data[5]~69 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[5]~70 (
	.dataa(\cmd_data[5]~69_combout ),
	.datab(csr_rd_inst_data_5),
	.datac(\cmd_data[2]~33_combout ),
	.datad(\cmd_data[2]~34_combout ),
	.cin(gnd),
	.combout(\cmd_data[5]~70_combout ),
	.cout());
defparam \cmd_data[5]~70 .lut_mask = 16'hCFA0;
defparam \cmd_data[5]~70 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[6]~72 (
	.dataa(csr_wr_inst_data_6),
	.datab(current_stateSTATE_WR_CMD),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\cmd_data[6]~72_combout ),
	.cout());
defparam \cmd_data[6]~72 .lut_mask = 16'h8888;
defparam \cmd_data[6]~72 .sum_lutc_input = "datac";

dffeas \mem_write_data_reg[6] (
	.clk(clk_clk),
	.d(avl_mem_writedata_6),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(\mem_write_data_reg[6]~q ),
	.prn(vcc));
defparam \mem_write_data_reg[6] .is_wysiwyg = "true";
defparam \mem_write_data_reg[6] .power_up = "low";

cycloneive_lcell_comb \cmd_data[6]~73 (
	.dataa(mem_write_data_reg_22),
	.datab(\mem_write_data_reg[6]~q ),
	.datac(\cmd_data[2]~26_combout ),
	.datad(\cmd_data[2]~25_combout ),
	.cin(gnd),
	.combout(\cmd_data[6]~73_combout ),
	.cout());
defparam \cmd_data[6]~73 .lut_mask = 16'h0AFC;
defparam \cmd_data[6]~73 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[6]~74 (
	.dataa(gnd),
	.datab(\mem_write_data_reg[14]~q ),
	.datac(mem_byteenable_reg_2),
	.datad(gnd),
	.cin(gnd),
	.combout(\cmd_data[6]~74_combout ),
	.cout());
defparam \cmd_data[6]~74 .lut_mask = 16'h0C0C;
defparam \cmd_data[6]~74 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[6]~75 (
	.dataa(mem_write_data_reg_30),
	.datab(\cmd_data[2]~28_combout ),
	.datac(\cmd_data[6]~74_combout ),
	.datad(\cmd_data[6]~73_combout ),
	.cin(gnd),
	.combout(\cmd_data[6]~75_combout ),
	.cout());
defparam \cmd_data[6]~75 .lut_mask = 16'h0C88;
defparam \cmd_data[6]~75 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[6]~76 (
	.dataa(mem_byteenable_reg_0),
	.datab(\cmd_data[2]~25_combout ),
	.datac(\cmd_data[6]~73_combout ),
	.datad(\cmd_data[6]~75_combout ),
	.cin(gnd),
	.combout(\cmd_data[6]~76_combout ),
	.cout());
defparam \cmd_data[6]~76 .lut_mask = 16'h0570;
defparam \cmd_data[6]~76 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[6]~77 (
	.dataa(\cmd_data[6]~76_combout ),
	.datab(csr_rd_inst_data_6),
	.datac(\cmd_data[2]~33_combout ),
	.datad(\cmd_data[2]~34_combout ),
	.cin(gnd),
	.combout(\cmd_data[6]~77_combout ),
	.cout());
defparam \cmd_data[6]~77 .lut_mask = 16'hCFA0;
defparam \cmd_data[6]~77 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[7]~79 (
	.dataa(csr_wr_inst_data_7),
	.datab(current_stateSTATE_WR_CMD),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\cmd_data[7]~79_combout ),
	.cout());
defparam \cmd_data[7]~79 .lut_mask = 16'h8888;
defparam \cmd_data[7]~79 .sum_lutc_input = "datac";

dffeas \mem_write_data_reg[7] (
	.clk(clk_clk),
	.d(avl_mem_writedata_7),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_wr_combi~0_combout ),
	.q(\mem_write_data_reg[7]~q ),
	.prn(vcc));
defparam \mem_write_data_reg[7] .is_wysiwyg = "true";
defparam \mem_write_data_reg[7] .power_up = "low";

cycloneive_lcell_comb \cmd_data[7]~80 (
	.dataa(mem_write_data_reg_23),
	.datab(\mem_write_data_reg[7]~q ),
	.datac(\cmd_data[2]~26_combout ),
	.datad(\cmd_data[2]~25_combout ),
	.cin(gnd),
	.combout(\cmd_data[7]~80_combout ),
	.cout());
defparam \cmd_data[7]~80 .lut_mask = 16'h0AFC;
defparam \cmd_data[7]~80 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[7]~81 (
	.dataa(gnd),
	.datab(\mem_write_data_reg[15]~q ),
	.datac(mem_byteenable_reg_2),
	.datad(gnd),
	.cin(gnd),
	.combout(\cmd_data[7]~81_combout ),
	.cout());
defparam \cmd_data[7]~81 .lut_mask = 16'h0C0C;
defparam \cmd_data[7]~81 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[7]~82 (
	.dataa(mem_write_data_reg_31),
	.datab(\cmd_data[2]~28_combout ),
	.datac(\cmd_data[7]~81_combout ),
	.datad(\cmd_data[7]~80_combout ),
	.cin(gnd),
	.combout(\cmd_data[7]~82_combout ),
	.cout());
defparam \cmd_data[7]~82 .lut_mask = 16'h0C88;
defparam \cmd_data[7]~82 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[7]~83 (
	.dataa(mem_byteenable_reg_0),
	.datab(\cmd_data[2]~25_combout ),
	.datac(\cmd_data[7]~80_combout ),
	.datad(\cmd_data[7]~82_combout ),
	.cin(gnd),
	.combout(\cmd_data[7]~83_combout ),
	.cout());
defparam \cmd_data[7]~83 .lut_mask = 16'h0570;
defparam \cmd_data[7]~83 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[7]~84 (
	.dataa(\cmd_data[7]~83_combout ),
	.datab(csr_rd_inst_data_7),
	.datac(\cmd_data[2]~33_combout ),
	.datad(\cmd_data[2]~34_combout ),
	.cin(gnd),
	.combout(\cmd_data[7]~84_combout ),
	.cout());
defparam \cmd_data[7]~84 .lut_mask = 16'hCFA0;
defparam \cmd_data[7]~84 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[12]~86 (
	.dataa(mem_byteenable_reg_3),
	.datab(mem_byteenable_reg_2),
	.datac(mem_write_data_reg_28),
	.datad(mem_byteenable_reg_0),
	.cin(gnd),
	.combout(\cmd_data[12]~86_combout ),
	.cout());
defparam \cmd_data[12]~86 .lut_mask = 16'h0080;
defparam \cmd_data[12]~86 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector16~0 (
	.dataa(csr_rd_inst_data_9),
	.datab(csr_rd_inst_data_10),
	.datac(csr_rd_inst_data_11),
	.datad(csr_rd_inst_data_12),
	.cin(gnd),
	.combout(\Selector16~0_combout ),
	.cout());
defparam \Selector16~0 .lut_mask = 16'hFFFE;
defparam \Selector16~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector16~1 (
	.dataa(current_stateSTATE_READ_CMD),
	.datab(csr_rd_inst_data_8),
	.datac(\Selector16~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector16~1_combout ),
	.cout());
defparam \Selector16~1 .lut_mask = 16'hA8A8;
defparam \Selector16~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \cmd_data[12]~87 (
	.dataa(\Selector16~1_combout ),
	.datab(\avst_fifo_inst|avst_fifo|out_payload[12]~q ),
	.datac(\cmd_data[8]~6_combout ),
	.datad(\cmd_data[8]~5_combout ),
	.cin(gnd),
	.combout(\cmd_data[12]~87_combout ),
	.cout());
defparam \cmd_data[12]~87 .lut_mask = 16'hA0CF;
defparam \cmd_data[12]~87 .sum_lutc_input = "datac";

endmodule

module flashLoader_avst_fifo (
	altera_reset_synchronizer_int_chain_out,
	Equal2,
	full,
	saved_grant_0,
	out_valid,
	current_stateSTATE_WR_DATA,
	Selector18,
	adap_out_cmd_ready,
	Selector181,
	mem_wr_combi,
	sink0_ready,
	out_payload_30,
	out_payload_29,
	out_payload_28,
	out_payload_27,
	out_payload_32,
	fifo_in_valid,
	out_payload_11,
	out_payload_18,
	out_payload_19,
	out_payload_21,
	out_payload_20,
	out_payload_22,
	out_payload_23,
	out_payload_24,
	out_payload_25,
	out_payload_26,
	out_payload_10,
	out_payload_8,
	out_payload_13,
	out_payload_17,
	out_payload_16,
	out_payload_15,
	out_payload_14,
	out_payload_9,
	out_payload_0,
	out_payload_4,
	out_payload_2,
	out_payload_1,
	out_payload_3,
	out_payload_5,
	out_payload_6,
	out_payload_7,
	out_payload_12,
	out_payload_31,
	clk_clk,
	avl_mem_writedata_30,
	avl_mem_writedata_29,
	avl_mem_writedata_28,
	avl_mem_writedata_27,
	avl_mem_writedata_11,
	avl_mem_writedata_18,
	avl_mem_writedata_19,
	avl_mem_writedata_21,
	avl_mem_writedata_20,
	avl_mem_writedata_22,
	avl_mem_writedata_23,
	avl_mem_writedata_24,
	avl_mem_writedata_25,
	avl_mem_writedata_26,
	avl_mem_writedata_10,
	avl_mem_writedata_8,
	avl_mem_writedata_13,
	avl_mem_writedata_17,
	avl_mem_writedata_16,
	avl_mem_writedata_15,
	avl_mem_writedata_31,
	avl_mem_writedata_14,
	avl_mem_writedata_9,
	avl_mem_writedata_0,
	avl_mem_writedata_4,
	avl_mem_writedata_12,
	avl_mem_writedata_2,
	avl_mem_writedata_1,
	avl_mem_writedata_3,
	avl_mem_writedata_5,
	avl_mem_writedata_6,
	avl_mem_writedata_7)/* synthesis synthesis_greybox=0 */;
input 	altera_reset_synchronizer_int_chain_out;
input 	Equal2;
output 	full;
input 	saved_grant_0;
output 	out_valid;
input 	current_stateSTATE_WR_DATA;
input 	Selector18;
input 	adap_out_cmd_ready;
input 	Selector181;
input 	mem_wr_combi;
input 	sink0_ready;
output 	out_payload_30;
output 	out_payload_29;
output 	out_payload_28;
output 	out_payload_27;
output 	out_payload_32;
input 	fifo_in_valid;
output 	out_payload_11;
output 	out_payload_18;
output 	out_payload_19;
output 	out_payload_21;
output 	out_payload_20;
output 	out_payload_22;
output 	out_payload_23;
output 	out_payload_24;
output 	out_payload_25;
output 	out_payload_26;
output 	out_payload_10;
output 	out_payload_8;
output 	out_payload_13;
output 	out_payload_17;
output 	out_payload_16;
output 	out_payload_15;
output 	out_payload_14;
output 	out_payload_9;
output 	out_payload_0;
output 	out_payload_4;
output 	out_payload_2;
output 	out_payload_1;
output 	out_payload_3;
output 	out_payload_5;
output 	out_payload_6;
output 	out_payload_7;
output 	out_payload_12;
output 	out_payload_31;
input 	clk_clk;
input 	avl_mem_writedata_30;
input 	avl_mem_writedata_29;
input 	avl_mem_writedata_28;
input 	avl_mem_writedata_27;
input 	avl_mem_writedata_11;
input 	avl_mem_writedata_18;
input 	avl_mem_writedata_19;
input 	avl_mem_writedata_21;
input 	avl_mem_writedata_20;
input 	avl_mem_writedata_22;
input 	avl_mem_writedata_23;
input 	avl_mem_writedata_24;
input 	avl_mem_writedata_25;
input 	avl_mem_writedata_26;
input 	avl_mem_writedata_10;
input 	avl_mem_writedata_8;
input 	avl_mem_writedata_13;
input 	avl_mem_writedata_17;
input 	avl_mem_writedata_16;
input 	avl_mem_writedata_15;
input 	avl_mem_writedata_31;
input 	avl_mem_writedata_14;
input 	avl_mem_writedata_9;
input 	avl_mem_writedata_0;
input 	avl_mem_writedata_4;
input 	avl_mem_writedata_12;
input 	avl_mem_writedata_2;
input 	avl_mem_writedata_1;
input 	avl_mem_writedata_3;
input 	avl_mem_writedata_5;
input 	avl_mem_writedata_6;
input 	avl_mem_writedata_7;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



flashLoader_altera_avalon_sc_fifo_1 avst_fifo(
	.reset(altera_reset_synchronizer_int_chain_out),
	.Equal2(Equal2),
	.full1(full),
	.saved_grant_0(saved_grant_0),
	.out_valid1(out_valid),
	.current_stateSTATE_WR_DATA(current_stateSTATE_WR_DATA),
	.Selector18(Selector18),
	.adap_out_cmd_ready(adap_out_cmd_ready),
	.Selector181(Selector181),
	.mem_wr_combi(mem_wr_combi),
	.sink0_ready(sink0_ready),
	.out_payload_30(out_payload_30),
	.out_payload_29(out_payload_29),
	.out_payload_28(out_payload_28),
	.out_payload_27(out_payload_27),
	.out_payload_32(out_payload_32),
	.fifo_in_valid(fifo_in_valid),
	.out_payload_11(out_payload_11),
	.out_payload_18(out_payload_18),
	.out_payload_19(out_payload_19),
	.out_payload_21(out_payload_21),
	.out_payload_20(out_payload_20),
	.out_payload_22(out_payload_22),
	.out_payload_23(out_payload_23),
	.out_payload_24(out_payload_24),
	.out_payload_25(out_payload_25),
	.out_payload_26(out_payload_26),
	.out_payload_10(out_payload_10),
	.out_payload_8(out_payload_8),
	.out_payload_13(out_payload_13),
	.out_payload_17(out_payload_17),
	.out_payload_16(out_payload_16),
	.out_payload_15(out_payload_15),
	.out_payload_14(out_payload_14),
	.out_payload_9(out_payload_9),
	.out_payload_0(out_payload_0),
	.out_payload_4(out_payload_4),
	.out_payload_2(out_payload_2),
	.out_payload_1(out_payload_1),
	.out_payload_3(out_payload_3),
	.out_payload_5(out_payload_5),
	.out_payload_6(out_payload_6),
	.out_payload_7(out_payload_7),
	.out_payload_12(out_payload_12),
	.out_payload_31(out_payload_31),
	.clk(clk_clk),
	.avl_mem_writedata_30(avl_mem_writedata_30),
	.avl_mem_writedata_29(avl_mem_writedata_29),
	.avl_mem_writedata_28(avl_mem_writedata_28),
	.avl_mem_writedata_27(avl_mem_writedata_27),
	.avl_mem_writedata_11(avl_mem_writedata_11),
	.avl_mem_writedata_18(avl_mem_writedata_18),
	.avl_mem_writedata_19(avl_mem_writedata_19),
	.avl_mem_writedata_21(avl_mem_writedata_21),
	.avl_mem_writedata_20(avl_mem_writedata_20),
	.avl_mem_writedata_22(avl_mem_writedata_22),
	.avl_mem_writedata_23(avl_mem_writedata_23),
	.avl_mem_writedata_24(avl_mem_writedata_24),
	.avl_mem_writedata_25(avl_mem_writedata_25),
	.avl_mem_writedata_26(avl_mem_writedata_26),
	.avl_mem_writedata_10(avl_mem_writedata_10),
	.avl_mem_writedata_8(avl_mem_writedata_8),
	.avl_mem_writedata_13(avl_mem_writedata_13),
	.avl_mem_writedata_17(avl_mem_writedata_17),
	.avl_mem_writedata_16(avl_mem_writedata_16),
	.avl_mem_writedata_15(avl_mem_writedata_15),
	.avl_mem_writedata_31(avl_mem_writedata_31),
	.avl_mem_writedata_14(avl_mem_writedata_14),
	.avl_mem_writedata_9(avl_mem_writedata_9),
	.avl_mem_writedata_0(avl_mem_writedata_0),
	.avl_mem_writedata_4(avl_mem_writedata_4),
	.avl_mem_writedata_12(avl_mem_writedata_12),
	.avl_mem_writedata_2(avl_mem_writedata_2),
	.avl_mem_writedata_1(avl_mem_writedata_1),
	.avl_mem_writedata_3(avl_mem_writedata_3),
	.avl_mem_writedata_5(avl_mem_writedata_5),
	.avl_mem_writedata_6(avl_mem_writedata_6),
	.avl_mem_writedata_7(avl_mem_writedata_7));

endmodule

module flashLoader_altera_avalon_sc_fifo_1 (
	reset,
	Equal2,
	full1,
	saved_grant_0,
	out_valid1,
	current_stateSTATE_WR_DATA,
	Selector18,
	adap_out_cmd_ready,
	Selector181,
	mem_wr_combi,
	sink0_ready,
	out_payload_30,
	out_payload_29,
	out_payload_28,
	out_payload_27,
	out_payload_32,
	fifo_in_valid,
	out_payload_11,
	out_payload_18,
	out_payload_19,
	out_payload_21,
	out_payload_20,
	out_payload_22,
	out_payload_23,
	out_payload_24,
	out_payload_25,
	out_payload_26,
	out_payload_10,
	out_payload_8,
	out_payload_13,
	out_payload_17,
	out_payload_16,
	out_payload_15,
	out_payload_14,
	out_payload_9,
	out_payload_0,
	out_payload_4,
	out_payload_2,
	out_payload_1,
	out_payload_3,
	out_payload_5,
	out_payload_6,
	out_payload_7,
	out_payload_12,
	out_payload_31,
	clk,
	avl_mem_writedata_30,
	avl_mem_writedata_29,
	avl_mem_writedata_28,
	avl_mem_writedata_27,
	avl_mem_writedata_11,
	avl_mem_writedata_18,
	avl_mem_writedata_19,
	avl_mem_writedata_21,
	avl_mem_writedata_20,
	avl_mem_writedata_22,
	avl_mem_writedata_23,
	avl_mem_writedata_24,
	avl_mem_writedata_25,
	avl_mem_writedata_26,
	avl_mem_writedata_10,
	avl_mem_writedata_8,
	avl_mem_writedata_13,
	avl_mem_writedata_17,
	avl_mem_writedata_16,
	avl_mem_writedata_15,
	avl_mem_writedata_31,
	avl_mem_writedata_14,
	avl_mem_writedata_9,
	avl_mem_writedata_0,
	avl_mem_writedata_4,
	avl_mem_writedata_12,
	avl_mem_writedata_2,
	avl_mem_writedata_1,
	avl_mem_writedata_3,
	avl_mem_writedata_5,
	avl_mem_writedata_6,
	avl_mem_writedata_7)/* synthesis synthesis_greybox=0 */;
input 	reset;
input 	Equal2;
output 	full1;
input 	saved_grant_0;
output 	out_valid1;
input 	current_stateSTATE_WR_DATA;
input 	Selector18;
input 	adap_out_cmd_ready;
input 	Selector181;
input 	mem_wr_combi;
input 	sink0_ready;
output 	out_payload_30;
output 	out_payload_29;
output 	out_payload_28;
output 	out_payload_27;
output 	out_payload_32;
input 	fifo_in_valid;
output 	out_payload_11;
output 	out_payload_18;
output 	out_payload_19;
output 	out_payload_21;
output 	out_payload_20;
output 	out_payload_22;
output 	out_payload_23;
output 	out_payload_24;
output 	out_payload_25;
output 	out_payload_26;
output 	out_payload_10;
output 	out_payload_8;
output 	out_payload_13;
output 	out_payload_17;
output 	out_payload_16;
output 	out_payload_15;
output 	out_payload_14;
output 	out_payload_9;
output 	out_payload_0;
output 	out_payload_4;
output 	out_payload_2;
output 	out_payload_1;
output 	out_payload_3;
output 	out_payload_5;
output 	out_payload_6;
output 	out_payload_7;
output 	out_payload_12;
output 	out_payload_31;
input 	clk;
input 	avl_mem_writedata_30;
input 	avl_mem_writedata_29;
input 	avl_mem_writedata_28;
input 	avl_mem_writedata_27;
input 	avl_mem_writedata_11;
input 	avl_mem_writedata_18;
input 	avl_mem_writedata_19;
input 	avl_mem_writedata_21;
input 	avl_mem_writedata_20;
input 	avl_mem_writedata_22;
input 	avl_mem_writedata_23;
input 	avl_mem_writedata_24;
input 	avl_mem_writedata_25;
input 	avl_mem_writedata_26;
input 	avl_mem_writedata_10;
input 	avl_mem_writedata_8;
input 	avl_mem_writedata_13;
input 	avl_mem_writedata_17;
input 	avl_mem_writedata_16;
input 	avl_mem_writedata_15;
input 	avl_mem_writedata_31;
input 	avl_mem_writedata_14;
input 	avl_mem_writedata_9;
input 	avl_mem_writedata_0;
input 	avl_mem_writedata_4;
input 	avl_mem_writedata_12;
input 	avl_mem_writedata_2;
input 	avl_mem_writedata_1;
input 	avl_mem_writedata_3;
input 	avl_mem_writedata_5;
input 	avl_mem_writedata_6;
input 	avl_mem_writedata_7;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read~0_combout ;
wire \wr_ptr[0]~0_combout ;
wire \wr_ptr[0]~q ;
wire \Add0~5_combout ;
wire \wr_ptr[1]~q ;
wire \mem_rd_ptr[0]~2_combout ;
wire \mem_rd_ptr[0]~3_combout ;
wire \rd_ptr[0]~q ;
wire \mem_rd_ptr[1]~0_combout ;
wire \mem_rd_ptr[1]~1_combout ;
wire \rd_ptr[1]~q ;
wire \internal_out_valid~0_combout ;
wire \Add0~4_combout ;
wire \wr_ptr[2]~q ;
wire \Add0~2_combout ;
wire \wr_ptr[3]~q ;
wire \mem_rd_ptr[3]~6_combout ;
wire \mem_rd_ptr[3]~7_combout ;
wire \rd_ptr[3]~q ;
wire \mem_rd_ptr[2]~10_combout ;
wire \mem_rd_ptr[2]~11_combout ;
wire \rd_ptr[2]~q ;
wire \Add1~0_combout ;
wire \internal_out_valid~1_combout ;
wire \Add1~1_combout ;
wire \mem_rd_ptr[4]~4_combout ;
wire \mem_rd_ptr[4]~5_combout ;
wire \rd_ptr[4]~q ;
wire \mem_rd_ptr[5]~8_combout ;
wire \mem_rd_ptr[5]~9_combout ;
wire \rd_ptr[5]~q ;
wire \Add0~0_combout ;
wire \Add0~1_combout ;
wire \wr_ptr[4]~q ;
wire \Add0~3_combout ;
wire \wr_ptr[5]~q ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \Equal0~2_combout ;
wire \internal_out_valid~2_combout ;
wire \next_empty~0_combout ;
wire \empty~q ;
wire \internal_out_valid~3_combout ;
wire \internal_out_valid~4_combout ;
wire \internal_out_valid~q ;
wire \next_full~0_combout ;
wire \next_full~1_combout ;
wire \next_full~2_combout ;
wire \next_full~3_combout ;
wire \next_full~4_combout ;
wire \next_full~5_combout ;
wire \internal_out_ready~0_combout ;
wire \internal_out_ready~combout ;
wire \mem_rtl_0|auto_generated|ram_block1a30~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a29~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a28~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a27~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a32~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a11~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a18~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a19~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a21~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a20~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a22~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a23~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a24~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a25~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a26~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a10~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a8~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a13~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a17~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a16~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a15~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a14~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a9~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a0~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a4~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a2~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a1~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a3~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a5~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a6~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a7~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a12~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a31~portbdataout ;

wire [143:0] \mem_rtl_0|auto_generated|ram_block1a30_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a29_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a28_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a27_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a32_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a11_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a18_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a19_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a21_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a20_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a22_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a23_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a24_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a25_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a26_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a10_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a8_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a13_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a17_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a16_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a15_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a14_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a9_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a2_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a1_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a3_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a5_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a6_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a7_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a12_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a31_PORTBDATAOUT_bus ;

assign \mem_rtl_0|auto_generated|ram_block1a30~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a30_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a29~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a29_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a28~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a28_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a27~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a27_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a32~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a32_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a11~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a11_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a18~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a18_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a19~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a19_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a21~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a21_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a20~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a20_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a22~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a22_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a23~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a23_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a24~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a24_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a25~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a25_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a26~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a26_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a10~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a10_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a8~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a8_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a13~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a13_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a17~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a17_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a16~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a16_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a15~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a15_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a14~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a14_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a9~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a9_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a0~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a4~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a2~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a2_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a1~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a1_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a3~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a3_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a5~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a5_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a6~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a6_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a7~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a7_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a12~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a12_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a31~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a31_PORTBDATAOUT_bus [0];

dffeas full(
	.clk(clk),
	.d(\next_full~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(full1),
	.prn(vcc));
defparam full.is_wysiwyg = "true";
defparam full.power_up = "low";

dffeas out_valid(
	.clk(clk),
	.d(\internal_out_valid~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_valid1),
	.prn(vcc));
defparam out_valid.is_wysiwyg = "true";
defparam out_valid.power_up = "low";

dffeas \out_payload[30] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a30~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_30),
	.prn(vcc));
defparam \out_payload[30] .is_wysiwyg = "true";
defparam \out_payload[30] .power_up = "low";

dffeas \out_payload[29] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a29~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_29),
	.prn(vcc));
defparam \out_payload[29] .is_wysiwyg = "true";
defparam \out_payload[29] .power_up = "low";

dffeas \out_payload[28] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a28~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_28),
	.prn(vcc));
defparam \out_payload[28] .is_wysiwyg = "true";
defparam \out_payload[28] .power_up = "low";

dffeas \out_payload[27] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a27~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_27),
	.prn(vcc));
defparam \out_payload[27] .is_wysiwyg = "true";
defparam \out_payload[27] .power_up = "low";

dffeas \out_payload[32] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a32~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_32),
	.prn(vcc));
defparam \out_payload[32] .is_wysiwyg = "true";
defparam \out_payload[32] .power_up = "low";

dffeas \out_payload[11] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a11~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_11),
	.prn(vcc));
defparam \out_payload[11] .is_wysiwyg = "true";
defparam \out_payload[11] .power_up = "low";

dffeas \out_payload[18] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a18~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_18),
	.prn(vcc));
defparam \out_payload[18] .is_wysiwyg = "true";
defparam \out_payload[18] .power_up = "low";

dffeas \out_payload[19] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a19~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_19),
	.prn(vcc));
defparam \out_payload[19] .is_wysiwyg = "true";
defparam \out_payload[19] .power_up = "low";

dffeas \out_payload[21] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a21~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_21),
	.prn(vcc));
defparam \out_payload[21] .is_wysiwyg = "true";
defparam \out_payload[21] .power_up = "low";

dffeas \out_payload[20] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a20~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_20),
	.prn(vcc));
defparam \out_payload[20] .is_wysiwyg = "true";
defparam \out_payload[20] .power_up = "low";

dffeas \out_payload[22] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a22~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_22),
	.prn(vcc));
defparam \out_payload[22] .is_wysiwyg = "true";
defparam \out_payload[22] .power_up = "low";

dffeas \out_payload[23] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a23~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_23),
	.prn(vcc));
defparam \out_payload[23] .is_wysiwyg = "true";
defparam \out_payload[23] .power_up = "low";

dffeas \out_payload[24] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a24~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_24),
	.prn(vcc));
defparam \out_payload[24] .is_wysiwyg = "true";
defparam \out_payload[24] .power_up = "low";

dffeas \out_payload[25] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a25~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_25),
	.prn(vcc));
defparam \out_payload[25] .is_wysiwyg = "true";
defparam \out_payload[25] .power_up = "low";

dffeas \out_payload[26] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a26~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_26),
	.prn(vcc));
defparam \out_payload[26] .is_wysiwyg = "true";
defparam \out_payload[26] .power_up = "low";

dffeas \out_payload[10] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a10~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_10),
	.prn(vcc));
defparam \out_payload[10] .is_wysiwyg = "true";
defparam \out_payload[10] .power_up = "low";

dffeas \out_payload[8] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a8~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_8),
	.prn(vcc));
defparam \out_payload[8] .is_wysiwyg = "true";
defparam \out_payload[8] .power_up = "low";

dffeas \out_payload[13] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a13~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_13),
	.prn(vcc));
defparam \out_payload[13] .is_wysiwyg = "true";
defparam \out_payload[13] .power_up = "low";

dffeas \out_payload[17] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a17~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_17),
	.prn(vcc));
defparam \out_payload[17] .is_wysiwyg = "true";
defparam \out_payload[17] .power_up = "low";

dffeas \out_payload[16] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a16~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_16),
	.prn(vcc));
defparam \out_payload[16] .is_wysiwyg = "true";
defparam \out_payload[16] .power_up = "low";

dffeas \out_payload[15] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a15~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_15),
	.prn(vcc));
defparam \out_payload[15] .is_wysiwyg = "true";
defparam \out_payload[15] .power_up = "low";

dffeas \out_payload[14] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a14~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_14),
	.prn(vcc));
defparam \out_payload[14] .is_wysiwyg = "true";
defparam \out_payload[14] .power_up = "low";

dffeas \out_payload[9] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a9~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_9),
	.prn(vcc));
defparam \out_payload[9] .is_wysiwyg = "true";
defparam \out_payload[9] .power_up = "low";

dffeas \out_payload[0] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a0~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_0),
	.prn(vcc));
defparam \out_payload[0] .is_wysiwyg = "true";
defparam \out_payload[0] .power_up = "low";

dffeas \out_payload[4] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a4~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_4),
	.prn(vcc));
defparam \out_payload[4] .is_wysiwyg = "true";
defparam \out_payload[4] .power_up = "low";

dffeas \out_payload[2] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a2~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_2),
	.prn(vcc));
defparam \out_payload[2] .is_wysiwyg = "true";
defparam \out_payload[2] .power_up = "low";

dffeas \out_payload[1] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a1~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_1),
	.prn(vcc));
defparam \out_payload[1] .is_wysiwyg = "true";
defparam \out_payload[1] .power_up = "low";

dffeas \out_payload[3] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a3~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_3),
	.prn(vcc));
defparam \out_payload[3] .is_wysiwyg = "true";
defparam \out_payload[3] .power_up = "low";

dffeas \out_payload[5] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a5~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_5),
	.prn(vcc));
defparam \out_payload[5] .is_wysiwyg = "true";
defparam \out_payload[5] .power_up = "low";

dffeas \out_payload[6] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a6~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_6),
	.prn(vcc));
defparam \out_payload[6] .is_wysiwyg = "true";
defparam \out_payload[6] .power_up = "low";

dffeas \out_payload[7] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a7~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_7),
	.prn(vcc));
defparam \out_payload[7] .is_wysiwyg = "true";
defparam \out_payload[7] .power_up = "low";

dffeas \out_payload[12] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a12~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_12),
	.prn(vcc));
defparam \out_payload[12] .is_wysiwyg = "true";
defparam \out_payload[12] .power_up = "low";

dffeas \out_payload[31] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a31~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_31),
	.prn(vcc));
defparam \out_payload[31] .is_wysiwyg = "true";
defparam \out_payload[31] .power_up = "low";

cycloneive_lcell_comb \read~0 (
	.dataa(\internal_out_valid~q ),
	.datab(current_stateSTATE_WR_DATA),
	.datac(sink0_ready),
	.datad(out_valid1),
	.cin(gnd),
	.combout(\read~0_combout ),
	.cout());
defparam \read~0 .lut_mask = 16'h80AA;
defparam \read~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_ptr[0]~0 (
	.dataa(\wr_ptr[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_ptr[0]~0_combout ),
	.cout());
defparam \wr_ptr[0]~0 .lut_mask = 16'h5555;
defparam \wr_ptr[0]~0 .sum_lutc_input = "datac";

dffeas \wr_ptr[0] (
	.clk(clk),
	.d(\wr_ptr[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_in_valid),
	.q(\wr_ptr[0]~q ),
	.prn(vcc));
defparam \wr_ptr[0] .is_wysiwyg = "true";
defparam \wr_ptr[0] .power_up = "low";

cycloneive_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\wr_ptr[1]~q ),
	.datad(\wr_ptr[0]~q ),
	.cin(gnd),
	.combout(\Add0~5_combout ),
	.cout());
defparam \Add0~5 .lut_mask = 16'h0FF0;
defparam \Add0~5 .sum_lutc_input = "datac";

dffeas \wr_ptr[1] (
	.clk(clk),
	.d(\Add0~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_in_valid),
	.q(\wr_ptr[1]~q ),
	.prn(vcc));
defparam \wr_ptr[1] .is_wysiwyg = "true";
defparam \wr_ptr[1] .power_up = "low";

cycloneive_lcell_comb \mem_rd_ptr[0]~2 (
	.dataa(\internal_out_valid~q ),
	.datab(current_stateSTATE_WR_DATA),
	.datac(out_valid1),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_rd_ptr[0]~2_combout ),
	.cout());
defparam \mem_rd_ptr[0]~2 .lut_mask = 16'h8A8A;
defparam \mem_rd_ptr[0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_rd_ptr[0]~3 (
	.dataa(\rd_ptr[0]~q ),
	.datab(sink0_ready),
	.datac(out_valid1),
	.datad(\mem_rd_ptr[0]~2_combout ),
	.cin(gnd),
	.combout(\mem_rd_ptr[0]~3_combout ),
	.cout());
defparam \mem_rd_ptr[0]~3 .lut_mask = 16'h65AA;
defparam \mem_rd_ptr[0]~3 .sum_lutc_input = "datac";

dffeas \rd_ptr[0] (
	.clk(clk),
	.d(\mem_rd_ptr[0]~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ptr[0]~q ),
	.prn(vcc));
defparam \rd_ptr[0] .is_wysiwyg = "true";
defparam \rd_ptr[0] .power_up = "low";

cycloneive_lcell_comb \mem_rd_ptr[1]~0 (
	.dataa(\rd_ptr[0]~q ),
	.datab(\internal_out_valid~q ),
	.datac(current_stateSTATE_WR_DATA),
	.datad(out_valid1),
	.cin(gnd),
	.combout(\mem_rd_ptr[1]~0_combout ),
	.cout());
defparam \mem_rd_ptr[1]~0 .lut_mask = 16'h8088;
defparam \mem_rd_ptr[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_rd_ptr[1]~1 (
	.dataa(\rd_ptr[1]~q ),
	.datab(sink0_ready),
	.datac(out_valid1),
	.datad(\mem_rd_ptr[1]~0_combout ),
	.cin(gnd),
	.combout(\mem_rd_ptr[1]~1_combout ),
	.cout());
defparam \mem_rd_ptr[1]~1 .lut_mask = 16'h65AA;
defparam \mem_rd_ptr[1]~1 .sum_lutc_input = "datac";

dffeas \rd_ptr[1] (
	.clk(clk),
	.d(\mem_rd_ptr[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ptr[1]~q ),
	.prn(vcc));
defparam \rd_ptr[1] .is_wysiwyg = "true";
defparam \rd_ptr[1] .power_up = "low";

cycloneive_lcell_comb \internal_out_valid~0 (
	.dataa(\wr_ptr[1]~q ),
	.datab(\rd_ptr[1]~q ),
	.datac(\wr_ptr[0]~q ),
	.datad(\rd_ptr[0]~q ),
	.cin(gnd),
	.combout(\internal_out_valid~0_combout ),
	.cout());
defparam \internal_out_valid~0 .lut_mask = 16'h0690;
defparam \internal_out_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~4 (
	.dataa(gnd),
	.datab(\wr_ptr[2]~q ),
	.datac(\wr_ptr[1]~q ),
	.datad(\wr_ptr[0]~q ),
	.cin(gnd),
	.combout(\Add0~4_combout ),
	.cout());
defparam \Add0~4 .lut_mask = 16'h3CCC;
defparam \Add0~4 .sum_lutc_input = "datac";

dffeas \wr_ptr[2] (
	.clk(clk),
	.d(\Add0~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_in_valid),
	.q(\wr_ptr[2]~q ),
	.prn(vcc));
defparam \wr_ptr[2] .is_wysiwyg = "true";
defparam \wr_ptr[2] .power_up = "low";

cycloneive_lcell_comb \Add0~2 (
	.dataa(\wr_ptr[3]~q ),
	.datab(\wr_ptr[2]~q ),
	.datac(\wr_ptr[1]~q ),
	.datad(\wr_ptr[0]~q ),
	.cin(gnd),
	.combout(\Add0~2_combout ),
	.cout());
defparam \Add0~2 .lut_mask = 16'h6AAA;
defparam \Add0~2 .sum_lutc_input = "datac";

dffeas \wr_ptr[3] (
	.clk(clk),
	.d(\Add0~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_in_valid),
	.q(\wr_ptr[3]~q ),
	.prn(vcc));
defparam \wr_ptr[3] .is_wysiwyg = "true";
defparam \wr_ptr[3] .power_up = "low";

cycloneive_lcell_comb \mem_rd_ptr[3]~6 (
	.dataa(current_stateSTATE_WR_DATA),
	.datab(out_valid1),
	.datac(sink0_ready),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_rd_ptr[3]~6_combout ),
	.cout());
defparam \mem_rd_ptr[3]~6 .lut_mask = 16'h4C4C;
defparam \mem_rd_ptr[3]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_rd_ptr[3]~7 (
	.dataa(\internal_out_valid~q ),
	.datab(\Add1~0_combout ),
	.datac(\rd_ptr[3]~q ),
	.datad(\mem_rd_ptr[3]~6_combout ),
	.cin(gnd),
	.combout(\mem_rd_ptr[3]~7_combout ),
	.cout());
defparam \mem_rd_ptr[3]~7 .lut_mask = 16'hF0D8;
defparam \mem_rd_ptr[3]~7 .sum_lutc_input = "datac";

dffeas \rd_ptr[3] (
	.clk(clk),
	.d(\mem_rd_ptr[3]~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ptr[3]~q ),
	.prn(vcc));
defparam \rd_ptr[3] .is_wysiwyg = "true";
defparam \rd_ptr[3] .power_up = "low";

cycloneive_lcell_comb \mem_rd_ptr[2]~10 (
	.dataa(current_stateSTATE_WR_DATA),
	.datab(out_valid1),
	.datac(\rd_ptr[0]~q ),
	.datad(sink0_ready),
	.cin(gnd),
	.combout(\mem_rd_ptr[2]~10_combout ),
	.cout());
defparam \mem_rd_ptr[2]~10 .lut_mask = 16'hB030;
defparam \mem_rd_ptr[2]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_rd_ptr[2]~11 (
	.dataa(\rd_ptr[1]~q ),
	.datab(\internal_out_valid~q ),
	.datac(\rd_ptr[2]~q ),
	.datad(\mem_rd_ptr[2]~10_combout ),
	.cin(gnd),
	.combout(\mem_rd_ptr[2]~11_combout ),
	.cout());
defparam \mem_rd_ptr[2]~11 .lut_mask = 16'h78F0;
defparam \mem_rd_ptr[2]~11 .sum_lutc_input = "datac";

dffeas \rd_ptr[2] (
	.clk(clk),
	.d(\mem_rd_ptr[2]~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ptr[2]~q ),
	.prn(vcc));
defparam \rd_ptr[2] .is_wysiwyg = "true";
defparam \rd_ptr[2] .power_up = "low";

cycloneive_lcell_comb \Add1~0 (
	.dataa(\rd_ptr[3]~q ),
	.datab(\rd_ptr[2]~q ),
	.datac(\rd_ptr[0]~q ),
	.datad(\rd_ptr[1]~q ),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout());
defparam \Add1~0 .lut_mask = 16'h6AAA;
defparam \Add1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \internal_out_valid~1 (
	.dataa(\internal_out_valid~0_combout ),
	.datab(\wr_ptr[3]~q ),
	.datac(\Add1~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\internal_out_valid~1_combout ),
	.cout());
defparam \internal_out_valid~1 .lut_mask = 16'h8282;
defparam \internal_out_valid~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add1~1 (
	.dataa(\rd_ptr[2]~q ),
	.datab(\rd_ptr[3]~q ),
	.datac(\rd_ptr[0]~q ),
	.datad(\rd_ptr[1]~q ),
	.cin(gnd),
	.combout(\Add1~1_combout ),
	.cout());
defparam \Add1~1 .lut_mask = 16'h8000;
defparam \Add1~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_rd_ptr[4]~4 (
	.dataa(\Add1~1_combout ),
	.datab(\internal_out_valid~q ),
	.datac(current_stateSTATE_WR_DATA),
	.datad(out_valid1),
	.cin(gnd),
	.combout(\mem_rd_ptr[4]~4_combout ),
	.cout());
defparam \mem_rd_ptr[4]~4 .lut_mask = 16'h8088;
defparam \mem_rd_ptr[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_rd_ptr[4]~5 (
	.dataa(\rd_ptr[4]~q ),
	.datab(sink0_ready),
	.datac(out_valid1),
	.datad(\mem_rd_ptr[4]~4_combout ),
	.cin(gnd),
	.combout(\mem_rd_ptr[4]~5_combout ),
	.cout());
defparam \mem_rd_ptr[4]~5 .lut_mask = 16'h65AA;
defparam \mem_rd_ptr[4]~5 .sum_lutc_input = "datac";

dffeas \rd_ptr[4] (
	.clk(clk),
	.d(\mem_rd_ptr[4]~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ptr[4]~q ),
	.prn(vcc));
defparam \rd_ptr[4] .is_wysiwyg = "true";
defparam \rd_ptr[4] .power_up = "low";

cycloneive_lcell_comb \mem_rd_ptr[5]~8 (
	.dataa(current_stateSTATE_WR_DATA),
	.datab(out_valid1),
	.datac(\rd_ptr[4]~q ),
	.datad(sink0_ready),
	.cin(gnd),
	.combout(\mem_rd_ptr[5]~8_combout ),
	.cout());
defparam \mem_rd_ptr[5]~8 .lut_mask = 16'hB030;
defparam \mem_rd_ptr[5]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_rd_ptr[5]~9 (
	.dataa(\Add1~1_combout ),
	.datab(\internal_out_valid~q ),
	.datac(\rd_ptr[5]~q ),
	.datad(\mem_rd_ptr[5]~8_combout ),
	.cin(gnd),
	.combout(\mem_rd_ptr[5]~9_combout ),
	.cout());
defparam \mem_rd_ptr[5]~9 .lut_mask = 16'h78F0;
defparam \mem_rd_ptr[5]~9 .sum_lutc_input = "datac";

dffeas \rd_ptr[5] (
	.clk(clk),
	.d(\mem_rd_ptr[5]~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ptr[5]~q ),
	.prn(vcc));
defparam \rd_ptr[5] .is_wysiwyg = "true";
defparam \rd_ptr[5] .power_up = "low";

cycloneive_lcell_comb \Add0~0 (
	.dataa(\wr_ptr[3]~q ),
	.datab(\wr_ptr[2]~q ),
	.datac(\wr_ptr[1]~q ),
	.datad(\wr_ptr[0]~q ),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout());
defparam \Add0~0 .lut_mask = 16'h8000;
defparam \Add0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\wr_ptr[4]~q ),
	.datad(\Add0~0_combout ),
	.cin(gnd),
	.combout(\Add0~1_combout ),
	.cout());
defparam \Add0~1 .lut_mask = 16'h0FF0;
defparam \Add0~1 .sum_lutc_input = "datac";

dffeas \wr_ptr[4] (
	.clk(clk),
	.d(\Add0~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_in_valid),
	.q(\wr_ptr[4]~q ),
	.prn(vcc));
defparam \wr_ptr[4] .is_wysiwyg = "true";
defparam \wr_ptr[4] .power_up = "low";

cycloneive_lcell_comb \Add0~3 (
	.dataa(gnd),
	.datab(\wr_ptr[5]~q ),
	.datac(\wr_ptr[4]~q ),
	.datad(\Add0~0_combout ),
	.cin(gnd),
	.combout(\Add0~3_combout ),
	.cout());
defparam \Add0~3 .lut_mask = 16'h3CCC;
defparam \Add0~3 .sum_lutc_input = "datac";

dffeas \wr_ptr[5] (
	.clk(clk),
	.d(\Add0~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_in_valid),
	.q(\wr_ptr[5]~q ),
	.prn(vcc));
defparam \wr_ptr[5] .is_wysiwyg = "true";
defparam \wr_ptr[5] .power_up = "low";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(\rd_ptr[4]~q ),
	.datab(\Add1~1_combout ),
	.datac(\rd_ptr[5]~q ),
	.datad(\wr_ptr[5]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h8778;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~1 (
	.dataa(\rd_ptr[0]~q ),
	.datab(\rd_ptr[1]~q ),
	.datac(\wr_ptr[2]~q ),
	.datad(\rd_ptr[2]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h8778;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~2 (
	.dataa(\wr_ptr[4]~q ),
	.datab(\rd_ptr[4]~q ),
	.datac(\Add1~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'h9696;
defparam \Equal0~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \internal_out_valid~2 (
	.dataa(\internal_out_valid~1_combout ),
	.datab(\Equal0~0_combout ),
	.datac(\Equal0~1_combout ),
	.datad(\Equal0~2_combout ),
	.cin(gnd),
	.combout(\internal_out_valid~2_combout ),
	.cout());
defparam \internal_out_valid~2 .lut_mask = 16'h0002;
defparam \internal_out_valid~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_empty~0 (
	.dataa(\read~0_combout ),
	.datab(\internal_out_valid~2_combout ),
	.datac(fifo_in_valid),
	.datad(\empty~q ),
	.cin(gnd),
	.combout(\next_empty~0_combout ),
	.cout());
defparam \next_empty~0 .lut_mask = 16'hF750;
defparam \next_empty~0 .sum_lutc_input = "datac";

dffeas empty(
	.clk(clk),
	.d(\next_empty~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty~q ),
	.prn(vcc));
defparam empty.is_wysiwyg = "true";
defparam empty.power_up = "low";

cycloneive_lcell_comb \internal_out_valid~3 (
	.dataa(\internal_out_valid~2_combout ),
	.datab(\internal_out_valid~q ),
	.datac(current_stateSTATE_WR_DATA),
	.datad(out_valid1),
	.cin(gnd),
	.combout(\internal_out_valid~3_combout ),
	.cout());
defparam \internal_out_valid~3 .lut_mask = 16'h8088;
defparam \internal_out_valid~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \internal_out_valid~4 (
	.dataa(\empty~q ),
	.datab(sink0_ready),
	.datac(out_valid1),
	.datad(\internal_out_valid~3_combout ),
	.cin(gnd),
	.combout(\internal_out_valid~4_combout ),
	.cout());
defparam \internal_out_valid~4 .lut_mask = 16'h20AA;
defparam \internal_out_valid~4 .sum_lutc_input = "datac";

dffeas internal_out_valid(
	.clk(clk),
	.d(\internal_out_valid~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_valid~q ),
	.prn(vcc));
defparam internal_out_valid.is_wysiwyg = "true";
defparam internal_out_valid.power_up = "low";

cycloneive_lcell_comb \next_full~0 (
	.dataa(\wr_ptr[1]~q ),
	.datab(\rd_ptr[1]~q ),
	.datac(\rd_ptr[0]~q ),
	.datad(\wr_ptr[0]~q ),
	.cin(gnd),
	.combout(\next_full~0_combout ),
	.cout());
defparam \next_full~0 .lut_mask = 16'h0690;
defparam \next_full~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_full~1 (
	.dataa(\rd_ptr[4]~q ),
	.datab(\Add0~1_combout ),
	.datac(\rd_ptr[3]~q ),
	.datad(\Add0~2_combout ),
	.cin(gnd),
	.combout(\next_full~1_combout ),
	.cout());
defparam \next_full~1 .lut_mask = 16'h9009;
defparam \next_full~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_full~2 (
	.dataa(\rd_ptr[5]~q ),
	.datab(\Add0~3_combout ),
	.datac(\rd_ptr[2]~q ),
	.datad(\Add0~4_combout ),
	.cin(gnd),
	.combout(\next_full~2_combout ),
	.cout());
defparam \next_full~2 .lut_mask = 16'h9009;
defparam \next_full~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_full~3 (
	.dataa(mem_wr_combi),
	.datab(\next_full~0_combout ),
	.datac(\next_full~1_combout ),
	.datad(\next_full~2_combout ),
	.cin(gnd),
	.combout(\next_full~3_combout ),
	.cout());
defparam \next_full~3 .lut_mask = 16'h8000;
defparam \next_full~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_full~4 (
	.dataa(full1),
	.datab(\internal_out_valid~q ),
	.datac(out_valid1),
	.datad(\next_full~3_combout ),
	.cin(gnd),
	.combout(\next_full~4_combout ),
	.cout());
defparam \next_full~4 .lut_mask = 16'hF3A2;
defparam \next_full~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \next_full~5 (
	.dataa(\internal_out_valid~q ),
	.datab(current_stateSTATE_WR_DATA),
	.datac(sink0_ready),
	.datad(\next_full~4_combout ),
	.cin(gnd),
	.combout(\next_full~5_combout ),
	.cout());
defparam \next_full~5 .lut_mask = 16'h7F00;
defparam \next_full~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \internal_out_ready~0 (
	.dataa(current_stateSTATE_WR_DATA),
	.datab(saved_grant_0),
	.datac(Selector18),
	.datad(Selector181),
	.cin(gnd),
	.combout(\internal_out_ready~0_combout ),
	.cout());
defparam \internal_out_ready~0 .lut_mask = 16'h8880;
defparam \internal_out_ready~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb internal_out_ready(
	.dataa(out_valid1),
	.datab(Selector18),
	.datac(adap_out_cmd_ready),
	.datad(\internal_out_ready~0_combout ),
	.cin(gnd),
	.combout(\internal_out_ready~combout ),
	.cout());
defparam internal_out_ready.lut_mask = 16'hFD55;
defparam internal_out_ready.sum_lutc_input = "datac";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a30 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_30}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a30_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a30 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a30 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a30 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a30 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a30 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a30 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a30 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a30 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a30 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a30 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a30 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a30 .port_a_first_bit_number = 30;
defparam \mem_rtl_0|auto_generated|ram_block1a30 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a30 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a30 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a30 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a30 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a30 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a30 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a30 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a30 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a30 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a30 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a30 .port_b_first_bit_number = 30;
defparam \mem_rtl_0|auto_generated|ram_block1a30 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a30 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a30 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a30 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a30 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a30 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a29 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_29}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a29_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a29 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a29 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a29 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a29 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a29 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a29 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a29 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a29 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a29 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a29 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a29 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a29 .port_a_first_bit_number = 29;
defparam \mem_rtl_0|auto_generated|ram_block1a29 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a29 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a29 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a29 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a29 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a29 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a29 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a29 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a29 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a29 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a29 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a29 .port_b_first_bit_number = 29;
defparam \mem_rtl_0|auto_generated|ram_block1a29 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a29 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a29 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a29 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a29 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a29 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a28 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_28}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a28_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a28 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a28 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a28 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a28 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a28 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a28 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a28 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a28 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a28 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a28 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a28 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a28 .port_a_first_bit_number = 28;
defparam \mem_rtl_0|auto_generated|ram_block1a28 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a28 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a28 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a28 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a28 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a28 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a28 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a28 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a28 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a28 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a28 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a28 .port_b_first_bit_number = 28;
defparam \mem_rtl_0|auto_generated|ram_block1a28 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a28 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a28 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a28 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a28 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a28 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a27 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_27}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a27_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a27 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a27 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a27 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a27 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a27 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a27 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a27 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a27 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a27 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a27 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a27 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a27 .port_a_first_bit_number = 27;
defparam \mem_rtl_0|auto_generated|ram_block1a27 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a27 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a27 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a27 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a27 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a27 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a27 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a27 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a27 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a27 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a27 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a27 .port_b_first_bit_number = 27;
defparam \mem_rtl_0|auto_generated|ram_block1a27 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a27 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a27 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a27 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a27 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a27 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a32 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Equal2}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a32_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a32 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a32 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a32 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a32 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a32 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a32 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a32 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a32 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a32 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a32 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a32 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a32 .port_a_first_bit_number = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a32 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a32 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a32 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a32 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a32 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a32 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a32 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a32 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a32 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a32 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a32 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a32 .port_b_first_bit_number = 32;
defparam \mem_rtl_0|auto_generated|ram_block1a32 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a32 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a32 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a32 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a32 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a32 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a11 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_11}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a11_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a11 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_first_bit_number = 11;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_first_bit_number = 11;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a11 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a18 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_18}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a18_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a18 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_a_first_bit_number = 18;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_first_bit_number = 18;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a18 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a19 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_19}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a19_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a19 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_a_first_bit_number = 19;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_first_bit_number = 19;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a19 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a21 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_21}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a21_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a21 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a21 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a21 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a21 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a21 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a21 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a21 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a21 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a21 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a21 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a21 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a21 .port_a_first_bit_number = 21;
defparam \mem_rtl_0|auto_generated|ram_block1a21 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a21 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a21 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a21 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a21 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a21 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a21 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a21 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a21 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a21 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a21 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a21 .port_b_first_bit_number = 21;
defparam \mem_rtl_0|auto_generated|ram_block1a21 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a21 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a21 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a21 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a21 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a21 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a20 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_20}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a20_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a20 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a20 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a20 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a20 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a20 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a20 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a20 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a20 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a20 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a20 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a20 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a20 .port_a_first_bit_number = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a20 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a20 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a20 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a20 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a20 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a20 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a20 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a20 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a20 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a20 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a20 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a20 .port_b_first_bit_number = 20;
defparam \mem_rtl_0|auto_generated|ram_block1a20 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a20 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a20 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a20 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a20 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a20 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a22 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_22}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a22_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a22 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a22 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a22 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a22 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a22 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a22 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a22 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a22 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a22 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a22 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a22 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a22 .port_a_first_bit_number = 22;
defparam \mem_rtl_0|auto_generated|ram_block1a22 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a22 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a22 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a22 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a22 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a22 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a22 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a22 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a22 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a22 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a22 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a22 .port_b_first_bit_number = 22;
defparam \mem_rtl_0|auto_generated|ram_block1a22 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a22 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a22 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a22 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a22 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a22 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a23 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_23}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a23_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a23 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a23 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a23 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a23 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a23 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a23 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a23 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a23 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a23 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a23 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a23 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a23 .port_a_first_bit_number = 23;
defparam \mem_rtl_0|auto_generated|ram_block1a23 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a23 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a23 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a23 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a23 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a23 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a23 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a23 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a23 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a23 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a23 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a23 .port_b_first_bit_number = 23;
defparam \mem_rtl_0|auto_generated|ram_block1a23 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a23 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a23 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a23 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a23 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a23 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a24 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_24}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a24_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a24 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a24 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a24 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a24 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a24 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a24 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a24 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a24 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a24 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a24 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a24 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a24 .port_a_first_bit_number = 24;
defparam \mem_rtl_0|auto_generated|ram_block1a24 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a24 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a24 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a24 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a24 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a24 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a24 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a24 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a24 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a24 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a24 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a24 .port_b_first_bit_number = 24;
defparam \mem_rtl_0|auto_generated|ram_block1a24 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a24 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a24 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a24 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a24 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a24 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a25 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_25}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a25_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a25 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a25 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a25 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a25 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a25 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a25 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a25 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a25 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a25 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a25 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a25 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a25 .port_a_first_bit_number = 25;
defparam \mem_rtl_0|auto_generated|ram_block1a25 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a25 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a25 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a25 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a25 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a25 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a25 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a25 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a25 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a25 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a25 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a25 .port_b_first_bit_number = 25;
defparam \mem_rtl_0|auto_generated|ram_block1a25 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a25 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a25 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a25 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a25 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a25 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a26 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_26}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a26_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a26 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a26 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a26 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a26 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a26 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a26 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a26 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a26 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a26 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a26 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a26 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a26 .port_a_first_bit_number = 26;
defparam \mem_rtl_0|auto_generated|ram_block1a26 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a26 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a26 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a26 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a26 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a26 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a26 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a26 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a26 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a26 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a26 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a26 .port_b_first_bit_number = 26;
defparam \mem_rtl_0|auto_generated|ram_block1a26 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a26 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a26 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a26 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a26 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a26 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a10 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_10}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a10_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a10 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_first_bit_number = 10;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_first_bit_number = 10;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a10 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a8 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_8}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a8_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a8 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_first_bit_number = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_first_bit_number = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a8 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a13 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_13}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a13_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a13 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_first_bit_number = 13;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_first_bit_number = 13;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a13 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a17 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_17}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a17_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a17 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_a_first_bit_number = 17;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_first_bit_number = 17;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a17 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a16 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_16}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a16_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a16 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_a_first_bit_number = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_first_bit_number = 16;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a16 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a15 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_15}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a15_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a15 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_first_bit_number = 15;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_first_bit_number = 15;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a15 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a14 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_14}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a14_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a14 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_first_bit_number = 14;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_first_bit_number = 14;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a14 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a9 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_9}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a9_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a9 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_first_bit_number = 9;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_first_bit_number = 9;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a9 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a0 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_0}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a0 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_first_bit_number = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_first_bit_number = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a4 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_4}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a4 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_first_bit_number = 4;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_first_bit_number = 4;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a2 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_2}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a2_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a2 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_first_bit_number = 2;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_first_bit_number = 2;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a1 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_1}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a1_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a1 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_first_bit_number = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_first_bit_number = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a3 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_3}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a3_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a3 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_first_bit_number = 3;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_first_bit_number = 3;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a5 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_5}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a5_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a5 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_first_bit_number = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_first_bit_number = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a6 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_6}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a6_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a6 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_first_bit_number = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_first_bit_number = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a7 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_7}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a7_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a7 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_first_bit_number = 7;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_first_bit_number = 7;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a12 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_12}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a12_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a12 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_first_bit_number = 12;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_first_bit_number = 12;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a12 .ram_block_type = "auto";

cycloneive_ram_block \mem_rtl_0|auto_generated|ram_block1a31 (
	.portawe(fifo_in_valid),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,avl_mem_writedata_31}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~9_combout ,\mem_rd_ptr[4]~5_combout ,\mem_rd_ptr[3]~7_combout ,\mem_rd_ptr[2]~11_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~3_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a31_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a31 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a31 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a31 .logical_ram_name = "flashLoader_intel_generic_serial_flash_interface_top_0:intel_generic_serial_flash_interface_top_0|flashLoader_intel_generic_serial_flash_interface_top_0_xip_controller:xip_controller|avst_fifo:avst_fifo_inst|altera_avalon_sc_fifo:avst_fifo|altsyncram:mem_rtl_0|altsyncram_ssg1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a31 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a31 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a31 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a31 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a31 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a31 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a31 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a31 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a31 .port_a_first_bit_number = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a31 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a31 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a31 .port_a_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a31 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a31 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a31 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a31 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a31 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a31 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a31 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a31 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a31 .port_b_first_bit_number = 31;
defparam \mem_rtl_0|auto_generated|ram_block1a31 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a31 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a31 .port_b_logical_ram_width = 33;
defparam \mem_rtl_0|auto_generated|ram_block1a31 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a31 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a31 .ram_block_type = "auto";

endmodule

module flashLoader_intel_generic_serial_flash_interface_cmd (
	data_num_lines_1,
	data_num_lines_2,
	addr_num_lines_2,
	addr_num_lines_1,
	csr_op_protocol_data_0,
	csr_flash_cmd_addr_data_0,
	reset,
	csr_op_protocol_data_1,
	csr_flash_cmd_addr_data_1,
	csr_flash_cmd_addr_data_2,
	csr_flash_cmd_addr_data_3,
	csr_flash_cmd_addr_data_4,
	csr_op_protocol_data_4,
	csr_op_protocol_data_5,
	csr_flash_cmd_addr_data_5,
	csr_flash_cmd_addr_data_6,
	csr_flash_cmd_addr_data_7,
	csr_op_protocol_data_8,
	csr_flash_cmd_addr_data_8,
	csr_flash_cmd_addr_data_9,
	csr_op_protocol_data_9,
	csr_flash_cmd_addr_data_10,
	csr_flash_cmd_addr_data_11,
	csr_op_protocol_data_12,
	csr_flash_cmd_addr_data_12,
	csr_flash_cmd_wr_data_0_data_12,
	csr_flash_cmd_wr_data_1_data_12,
	csr_flash_cmd_addr_data_13,
	csr_op_protocol_data_13,
	csr_flash_cmd_addr_data_14,
	csr_flash_cmd_addr_data_15,
	csr_op_protocol_data_16,
	csr_flash_cmd_addr_data_16,
	csr_flash_cmd_addr_data_17,
	csr_op_protocol_data_17,
	csr_flash_cmd_addr_data_18,
	csr_flash_cmd_addr_data_19,
	csr_flash_cmd_addr_data_20,
	csr_flash_cmd_addr_data_21,
	csr_flash_cmd_addr_data_22,
	csr_flash_cmd_addr_data_23,
	csr_flash_cmd_addr_data_24,
	csr_flash_cmd_addr_data_25,
	csr_flash_cmd_addr_data_26,
	csr_flash_cmd_addr_data_27,
	csr_flash_cmd_addr_data_28,
	csr_flash_cmd_addr_data_29,
	csr_flash_cmd_addr_data_30,
	csr_flash_cmd_addr_data_31,
	csr_flash_cmd_wr_data_0_data_31,
	csr_flash_cmd_wr_data_1_data_31,
	stateST_SEND_DUMMY_RSP,
	out_valid,
	out_endofpacket,
	in_cmd_channel_reg_1,
	stateST_WAIT_RSP,
	out_data_0,
	out_rsp_data_0,
	current_stateSTATE_READ_DATA,
	out_rsp_data_1,
	out_rsp_data_2,
	out_rsp_data_3,
	out_rsp_data_4,
	out_rsp_data_5,
	out_rsp_data_6,
	out_rsp_data_7,
	out_rsp_data_8,
	out_rsp_data_9,
	out_rsp_data_10,
	out_rsp_data_11,
	out_rsp_data_12,
	out_rsp_data_13,
	out_rsp_data_14,
	out_rsp_data_15,
	out_rsp_data_16,
	out_rsp_data_17,
	out_rsp_data_18,
	out_rsp_data_19,
	out_rsp_data_20,
	out_rsp_data_21,
	out_rsp_data_22,
	out_rsp_data_23,
	out_rsp_data_24,
	out_rsp_data_25,
	out_rsp_data_26,
	out_rsp_data_27,
	out_rsp_data_28,
	out_rsp_data_29,
	out_rsp_data_30,
	out_rsp_data_31,
	in_cmd_channel_reg_0,
	header_information_30,
	header_information_29,
	header_information_28,
	header_information_27,
	WideOr0,
	stateST_IDLE,
	in_cmd_channel,
	stateST_SEND_HEADER,
	current_stateSTATE_WR_CMD,
	current_stateSTATE_READ_CMD,
	src_startofpacket,
	src_valid,
	current_stateSTATE_WR_DATA,
	cmd_valid,
	stateST_SEND_DATA,
	stateST_SEND_ADDR,
	Selector18,
	op_num_lines_1,
	data_num_lines_0,
	op_num_lines_0,
	WideOr01,
	in_ready,
	op_num_lines_2,
	WideOr02,
	adap_out_cmd_ready,
	Selector181,
	stateST_SEND_DATA_1,
	stateST_SEND_DATA_0,
	Selector182,
	header_information_11,
	src_data_30,
	is_burst_reg,
	src_data_301,
	src_data_302,
	in_cmd_data,
	src_data_29,
	src_data_291,
	src_data_28,
	src_data_281,
	src_data_27,
	src_data_271,
	stateST_SEND_OPCODE,
	Selector8,
	demux_channel_2,
	sink_ready,
	addr_num_lines_0,
	WideOr03,
	out_rsp_valid,
	WideOr1,
	src_payload_0,
	WideOr04,
	WideOr05,
	WideOr06,
	out_rsp_data_01,
	out_rsp_data_110,
	out_rsp_data_210,
	out_rsp_data_32,
	out_rsp_data_41,
	out_rsp_data_51,
	out_rsp_data_61,
	out_rsp_data_71,
	header_information_13,
	header_information_17,
	header_information_16,
	header_information_15,
	header_information_14,
	src_data_11,
	cmd_data_11,
	src_data_19,
	src_data_191,
	src_data_21,
	src_data_211,
	src_data_20,
	src_data_201,
	WideOr07,
	src_data_10,
	cmd_data_10,
	has_addr,
	src_data_8,
	cmd_data_8,
	src_data_13,
	cmd_data_13,
	src_data_17,
	src_data_171,
	src_data_16,
	src_data_161,
	src_data_15,
	mem_write_data_reg_31,
	cmd_data_15,
	src_data_14,
	cmd_data_14,
	src_data_9,
	cmd_data_9,
	Selector20,
	Selector16,
	Selector12,
	Selector14,
	Selector15,
	Selector13,
	Selector11,
	Selector10,
	Selector9,
	Selector17,
	mem_addr_reg_6,
	mem_addr_reg_14,
	addr_bytes_xip_0,
	mem_addr_reg_10,
	mem_addr_reg_18,
	mem_addr_reg_2,
	mem_addr_reg_8,
	mem_addr_reg_16,
	mem_addr_reg_0,
	mem_addr_reg_15,
	mem_addr_reg_7,
	WideOr19,
	mem_addr_reg_17,
	mem_addr_reg_9,
	mem_addr_reg_1,
	mem_addr_reg_19,
	mem_addr_reg_11,
	mem_addr_reg_3,
	mem_addr_reg_12,
	mem_addr_reg_20,
	mem_addr_reg_4,
	mem_addr_reg_13,
	mem_addr_reg_5,
	has_dummy,
	cmd_data_12,
	out_payload_31,
	clk_clk)/* synthesis synthesis_greybox=0 */;
output 	data_num_lines_1;
output 	data_num_lines_2;
output 	addr_num_lines_2;
output 	addr_num_lines_1;
input 	csr_op_protocol_data_0;
input 	csr_flash_cmd_addr_data_0;
input 	reset;
input 	csr_op_protocol_data_1;
input 	csr_flash_cmd_addr_data_1;
input 	csr_flash_cmd_addr_data_2;
input 	csr_flash_cmd_addr_data_3;
input 	csr_flash_cmd_addr_data_4;
input 	csr_op_protocol_data_4;
input 	csr_op_protocol_data_5;
input 	csr_flash_cmd_addr_data_5;
input 	csr_flash_cmd_addr_data_6;
input 	csr_flash_cmd_addr_data_7;
input 	csr_op_protocol_data_8;
input 	csr_flash_cmd_addr_data_8;
input 	csr_flash_cmd_addr_data_9;
input 	csr_op_protocol_data_9;
input 	csr_flash_cmd_addr_data_10;
input 	csr_flash_cmd_addr_data_11;
input 	csr_op_protocol_data_12;
input 	csr_flash_cmd_addr_data_12;
input 	csr_flash_cmd_wr_data_0_data_12;
input 	csr_flash_cmd_wr_data_1_data_12;
input 	csr_flash_cmd_addr_data_13;
input 	csr_op_protocol_data_13;
input 	csr_flash_cmd_addr_data_14;
input 	csr_flash_cmd_addr_data_15;
input 	csr_op_protocol_data_16;
input 	csr_flash_cmd_addr_data_16;
input 	csr_flash_cmd_addr_data_17;
input 	csr_op_protocol_data_17;
input 	csr_flash_cmd_addr_data_18;
input 	csr_flash_cmd_addr_data_19;
input 	csr_flash_cmd_addr_data_20;
input 	csr_flash_cmd_addr_data_21;
input 	csr_flash_cmd_addr_data_22;
input 	csr_flash_cmd_addr_data_23;
input 	csr_flash_cmd_addr_data_24;
input 	csr_flash_cmd_addr_data_25;
input 	csr_flash_cmd_addr_data_26;
input 	csr_flash_cmd_addr_data_27;
input 	csr_flash_cmd_addr_data_28;
input 	csr_flash_cmd_addr_data_29;
input 	csr_flash_cmd_addr_data_30;
input 	csr_flash_cmd_addr_data_31;
input 	csr_flash_cmd_wr_data_0_data_31;
input 	csr_flash_cmd_wr_data_1_data_31;
output 	stateST_SEND_DUMMY_RSP;
output 	out_valid;
output 	out_endofpacket;
output 	in_cmd_channel_reg_1;
input 	stateST_WAIT_RSP;
output 	out_data_0;
output 	out_rsp_data_0;
input 	current_stateSTATE_READ_DATA;
output 	out_rsp_data_1;
output 	out_rsp_data_2;
output 	out_rsp_data_3;
output 	out_rsp_data_4;
output 	out_rsp_data_5;
output 	out_rsp_data_6;
output 	out_rsp_data_7;
output 	out_rsp_data_8;
output 	out_rsp_data_9;
output 	out_rsp_data_10;
output 	out_rsp_data_11;
output 	out_rsp_data_12;
output 	out_rsp_data_13;
output 	out_rsp_data_14;
output 	out_rsp_data_15;
output 	out_rsp_data_16;
output 	out_rsp_data_17;
output 	out_rsp_data_18;
output 	out_rsp_data_19;
output 	out_rsp_data_20;
output 	out_rsp_data_21;
output 	out_rsp_data_22;
output 	out_rsp_data_23;
output 	out_rsp_data_24;
output 	out_rsp_data_25;
output 	out_rsp_data_26;
output 	out_rsp_data_27;
output 	out_rsp_data_28;
output 	out_rsp_data_29;
output 	out_rsp_data_30;
output 	out_rsp_data_31;
output 	in_cmd_channel_reg_0;
output 	header_information_30;
output 	header_information_29;
output 	header_information_28;
output 	header_information_27;
input 	WideOr0;
output 	stateST_IDLE;
input 	[1:0] in_cmd_channel;
input 	stateST_SEND_HEADER;
input 	current_stateSTATE_WR_CMD;
input 	current_stateSTATE_READ_CMD;
input 	src_startofpacket;
input 	src_valid;
input 	current_stateSTATE_WR_DATA;
input 	cmd_valid;
output 	stateST_SEND_DATA;
output 	stateST_SEND_ADDR;
output 	Selector18;
output 	op_num_lines_1;
output 	data_num_lines_0;
output 	op_num_lines_0;
input 	WideOr01;
input 	in_ready;
output 	op_num_lines_2;
input 	WideOr02;
output 	adap_out_cmd_ready;
output 	Selector181;
input 	stateST_SEND_DATA_1;
input 	stateST_SEND_DATA_0;
output 	Selector182;
output 	header_information_11;
input 	src_data_30;
input 	is_burst_reg;
input 	src_data_301;
input 	src_data_302;
input 	[31:0] in_cmd_data;
input 	src_data_29;
input 	src_data_291;
input 	src_data_28;
input 	src_data_281;
input 	src_data_27;
input 	src_data_271;
output 	stateST_SEND_OPCODE;
output 	Selector8;
input 	demux_channel_2;
input 	sink_ready;
output 	addr_num_lines_0;
input 	WideOr03;
input 	out_rsp_valid;
input 	WideOr1;
input 	src_payload_0;
input 	WideOr04;
input 	WideOr05;
input 	WideOr06;
input 	out_rsp_data_01;
input 	out_rsp_data_110;
input 	out_rsp_data_210;
input 	out_rsp_data_32;
input 	out_rsp_data_41;
input 	out_rsp_data_51;
input 	out_rsp_data_61;
input 	out_rsp_data_71;
output 	header_information_13;
output 	header_information_17;
output 	header_information_16;
output 	header_information_15;
output 	header_information_14;
input 	src_data_11;
input 	cmd_data_11;
input 	src_data_19;
input 	src_data_191;
input 	src_data_21;
input 	src_data_211;
input 	src_data_20;
input 	src_data_201;
input 	WideOr07;
input 	src_data_10;
input 	cmd_data_10;
input 	has_addr;
input 	src_data_8;
input 	cmd_data_8;
input 	src_data_13;
input 	cmd_data_13;
input 	src_data_17;
input 	src_data_171;
input 	src_data_16;
input 	src_data_161;
input 	src_data_15;
input 	mem_write_data_reg_31;
input 	cmd_data_15;
input 	src_data_14;
input 	cmd_data_14;
input 	src_data_9;
input 	cmd_data_9;
output 	Selector20;
output 	Selector16;
output 	Selector12;
output 	Selector14;
output 	Selector15;
output 	Selector13;
output 	Selector11;
output 	Selector10;
output 	Selector9;
output 	Selector17;
input 	mem_addr_reg_6;
input 	mem_addr_reg_14;
input 	addr_bytes_xip_0;
input 	mem_addr_reg_10;
input 	mem_addr_reg_18;
input 	mem_addr_reg_2;
input 	mem_addr_reg_8;
input 	mem_addr_reg_16;
input 	mem_addr_reg_0;
input 	mem_addr_reg_15;
input 	mem_addr_reg_7;
input 	WideOr19;
input 	mem_addr_reg_17;
input 	mem_addr_reg_9;
input 	mem_addr_reg_1;
input 	mem_addr_reg_19;
input 	mem_addr_reg_11;
input 	mem_addr_reg_3;
input 	mem_addr_reg_12;
input 	mem_addr_reg_20;
input 	mem_addr_reg_4;
input 	mem_addr_reg_13;
input 	mem_addr_reg_5;
input 	has_dummy;
input 	cmd_data_12;
input 	out_payload_31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data_adapter_8_32_inst|out_data[1]~q ;
wire \data_adapter_8_32_inst|out_data[2]~q ;
wire \data_adapter_8_32_inst|out_data[3]~q ;
wire \data_adapter_8_32_inst|out_data[4]~q ;
wire \data_adapter_8_32_inst|out_data[5]~q ;
wire \data_adapter_8_32_inst|out_data[6]~q ;
wire \data_adapter_8_32_inst|out_data[7]~q ;
wire \data_adapter_8_32_inst|out_data[8]~q ;
wire \data_adapter_8_32_inst|out_data[9]~q ;
wire \data_adapter_8_32_inst|out_data[10]~q ;
wire \data_adapter_8_32_inst|out_data[11]~q ;
wire \data_adapter_8_32_inst|out_data[12]~q ;
wire \data_adapter_8_32_inst|out_data[13]~q ;
wire \data_adapter_8_32_inst|out_data[14]~q ;
wire \data_adapter_8_32_inst|out_data[15]~q ;
wire \data_adapter_8_32_inst|out_data[16]~q ;
wire \data_adapter_8_32_inst|out_data[17]~q ;
wire \data_adapter_8_32_inst|out_data[18]~q ;
wire \data_adapter_8_32_inst|out_data[19]~q ;
wire \data_adapter_8_32_inst|out_data[20]~q ;
wire \data_adapter_8_32_inst|out_data[21]~q ;
wire \data_adapter_8_32_inst|out_data[22]~q ;
wire \data_adapter_8_32_inst|out_data[23]~q ;
wire \data_adapter_8_32_inst|out_data[24]~q ;
wire \data_adapter_8_32_inst|out_data[25]~q ;
wire \data_adapter_8_32_inst|out_data[26]~q ;
wire \data_adapter_8_32_inst|out_data[27]~q ;
wire \data_adapter_8_32_inst|out_data[28]~q ;
wire \data_adapter_8_32_inst|out_data[29]~q ;
wire \data_adapter_8_32_inst|out_data[30]~q ;
wire \data_adapter_8_32_inst|out_data[31]~q ;
wire \data_adapter_8_32_inst|a_valid~q ;
wire \data_adapter_8_32_inst|a_ready~combout ;
wire \comb~0_combout ;
wire \data_adapter_32_8_inst|state_register[1]~q ;
wire \data_adapter_32_8_inst|state_register[0]~q ;
wire \data_adapter_32_8_inst|out_valid~q ;
wire \data_adapter_32_8_inst|a_valid~q ;
wire \comb~1_combout ;
wire \data_adapter_8_32_inst|in_ready~combout ;
wire \adap_in_cmd_valid~0_combout ;
wire \data_adapter_32_8_inst|out_data[0]~q ;
wire \data_adapter_32_8_inst|out_data[4]~q ;
wire \data_adapter_32_8_inst|out_data[2]~q ;
wire \data_adapter_32_8_inst|out_data[1]~q ;
wire \data_adapter_32_8_inst|out_data[3]~q ;
wire \data_adapter_32_8_inst|out_data[5]~q ;
wire \data_adapter_32_8_inst|out_data[6]~q ;
wire \data_adapter_32_8_inst|out_data[7]~q ;
wire \adap_in_cmd_data[8]~0_combout ;
wire \adap_in_cmd_data[16]~1_combout ;
wire \adap_in_cmd_data[0]~2_combout ;
wire \adap_in_cmd_data[24]~3_combout ;
wire \adap_in_cmd_data[12]~4_combout ;
wire \adap_in_cmd_data[12]~5_combout ;
wire \adap_in_cmd_data[12]~6_combout ;
wire \adap_in_cmd_data[20]~7_combout ;
wire \adap_in_cmd_data[4]~8_combout ;
wire \adap_in_cmd_data[28]~9_combout ;
wire \adap_in_cmd_data[10]~10_combout ;
wire \adap_in_cmd_data[18]~11_combout ;
wire \adap_in_cmd_data[2]~12_combout ;
wire \adap_in_cmd_data[26]~13_combout ;
wire \adap_in_cmd_data[17]~14_combout ;
wire \adap_in_cmd_data[9]~15_combout ;
wire \adap_in_cmd_data[1]~16_combout ;
wire \adap_in_cmd_data[25]~17_combout ;
wire \adap_in_cmd_data[19]~18_combout ;
wire \adap_in_cmd_data[11]~19_combout ;
wire \adap_in_cmd_data[3]~20_combout ;
wire \adap_in_cmd_data[27]~21_combout ;
wire \adap_in_cmd_data[21]~22_combout ;
wire \adap_in_cmd_data[13]~23_combout ;
wire \adap_in_cmd_data[5]~24_combout ;
wire \adap_in_cmd_data[29]~25_combout ;
wire \adap_in_cmd_data[14]~26_combout ;
wire \adap_in_cmd_data[22]~27_combout ;
wire \adap_in_cmd_data[6]~28_combout ;
wire \adap_in_cmd_data[30]~29_combout ;
wire \adap_in_cmd_data[23]~30_combout ;
wire \adap_in_cmd_data[15]~31_combout ;
wire \adap_in_cmd_data[7]~32_combout ;
wire \adap_in_cmd_data[31]~33_combout ;
wire \adap_in_cmd_data[31]~34_combout ;
wire \adap_in_cmd_data[31]~35_combout ;
wire \adap_in_cmd_data[31]~36_combout ;
wire \Equal12~0_combout ;
wire \Equal8~0_combout ;
wire \Equal5~0_combout ;
wire \data_num_lines[1]~0_combout ;
wire \Equal3~0_combout ;
wire \always2~0_combout ;
wire \always2~1_combout ;
wire \always0~0_combout ;
wire \always0~1_combout ;
wire \data_num_lines~7_combout ;
wire \data_num_lines~8_combout ;
wire \data_num_lines[2]~1_combout ;
wire \Equal4~0_combout ;
wire \addr_num_lines~4_combout ;
wire \addr_num_lines~5_combout ;
wire \addr_num_lines[2]~1_combout ;
wire \Equal10~0_combout ;
wire \Equal6~0_combout ;
wire \addr_num_lines[1]~0_combout ;
wire \header_information[18]~q ;
wire \Add2~0_combout ;
wire \header_information[19]~q ;
wire \Add2~1 ;
wire \Add2~2_combout ;
wire \data_in_cnt[0]~8_combout ;
wire \data_in_cnt_done~combout ;
wire \always8~0_combout ;
wire \data_in_cnt[0]~q ;
wire \data_in_cnt[0]~9 ;
wire \data_in_cnt[1]~10_combout ;
wire \data_in_cnt[1]~q ;
wire \data_in_cnt_done~0_combout ;
wire \header_information[21]~q ;
wire \header_information[20]~q ;
wire \Add2~3 ;
wire \Add2~5 ;
wire \Add2~6_combout ;
wire \data_in_cnt[1]~11 ;
wire \data_in_cnt[2]~12_combout ;
wire \data_in_cnt[2]~q ;
wire \data_in_cnt[2]~13 ;
wire \data_in_cnt[3]~14_combout ;
wire \data_in_cnt[3]~q ;
wire \Add2~4_combout ;
wire \Equal16~0_combout ;
wire \data_in_cnt_done~1_combout ;
wire \header_information[22]~q ;
wire \Add2~7 ;
wire \Add2~8_combout ;
wire \header_information[23]~q ;
wire \Add2~9 ;
wire \Add2~10_combout ;
wire \data_in_cnt[3]~15 ;
wire \data_in_cnt[4]~16_combout ;
wire \data_in_cnt[4]~q ;
wire \data_in_cnt[4]~17 ;
wire \data_in_cnt[5]~18_combout ;
wire \data_in_cnt[5]~q ;
wire \data_in_cnt_done~2_combout ;
wire \header_information[24]~q ;
wire \Add2~11 ;
wire \Add2~12_combout ;
wire \header_information[25]~q ;
wire \Add2~13 ;
wire \Add2~14_combout ;
wire \data_in_cnt[5]~19 ;
wire \data_in_cnt[6]~20_combout ;
wire \data_in_cnt[6]~q ;
wire \data_in_cnt[6]~21 ;
wire \data_in_cnt[7]~22_combout ;
wire \data_in_cnt[7]~q ;
wire \data_in_cnt_done~3_combout ;
wire \header_information[26]~q ;
wire \Add2~15 ;
wire \Add2~16_combout ;
wire \data_in_cnt_done~4_combout ;
wire \Selector5~2_combout ;
wire \Selector5~3_combout ;
wire \Selector5~7_combout ;
wire \Selector5~4_combout ;
wire \header_information[10]~q ;
wire \Selector5~5_combout ;
wire \header_information[8]~q ;
wire \Selector3~2_combout ;
wire \header_information[9]~q ;
wire \addr_cnt_done~0_combout ;
wire \addr_cnt_next[0]~1_combout ;
wire \addr_cnt_next[0]~2_combout ;
wire \addr_cnt[0]~q ;
wire \addr_cnt_next[1]~0_combout ;
wire \addr_cnt[1]~q ;
wire \Selector20~0_combout ;
wire \Selector20~1_combout ;
wire \Selector5~6_combout ;
wire \state.ST_WAIT_BUFFER~q ;
wire \buffer_cnt[0]~2_combout ;
wire \buffer_cnt[0]~q ;
wire \buffer_cnt[1]~1_combout ;
wire \buffer_cnt[1]~q ;
wire \buffer_cnt[2]~0_combout ;
wire \buffer_cnt[2]~q ;
wire \Selector6~0_combout ;
wire \Selector6~1_combout ;
wire \data_out_cnt[0]~8_combout ;
wire \always12~1_combout ;
wire \data_out_cnt[0]~q ;
wire \data_out_cnt[0]~9 ;
wire \data_out_cnt[1]~10_combout ;
wire \data_out_cnt[1]~q ;
wire \data_out_cnt[1]~11 ;
wire \data_out_cnt[2]~12_combout ;
wire \data_out_cnt[2]~q ;
wire \data_out_cnt[2]~13 ;
wire \data_out_cnt[3]~14_combout ;
wire \data_out_cnt[3]~q ;
wire \in_rsp_eop~0_combout ;
wire \data_out_cnt[3]~15 ;
wire \data_out_cnt[4]~16_combout ;
wire \data_out_cnt[4]~q ;
wire \data_out_cnt[4]~17 ;
wire \data_out_cnt[5]~18_combout ;
wire \data_out_cnt[5]~q ;
wire \data_out_cnt[5]~19 ;
wire \data_out_cnt[6]~20_combout ;
wire \data_out_cnt[6]~q ;
wire \in_rsp_eop~1_combout ;
wire \in_rsp_eop~2_combout ;
wire \data_out_cnt[6]~21 ;
wire \data_out_cnt[7]~22_combout ;
wire \data_out_cnt[7]~q ;
wire \in_rsp_eop~3_combout ;
wire \in_rsp_eop~4_combout ;
wire \in_rsp_eop~combout ;
wire \Selector4~0_combout ;
wire \Selector4~1_combout ;
wire \Selector4~2_combout ;
wire \state.ST_WAIT_RSP~q ;
wire \Selector7~0_combout ;
wire \Selector7~1_combout ;
wire \state.ST_COMPLETE~q ;
wire \Selector0~0_combout ;
wire \Selector0~1_combout ;
wire \Selector3~6_combout ;
wire \Selector3~3_combout ;
wire \Selector3~4_combout ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \Selector2~2_combout ;
wire \Selector18~0_combout ;
wire \last_word_detect~0_combout ;
wire \last_word_detect~1_combout ;
wire \last_word_detect~q ;
wire \Selector18~1_combout ;
wire \data_num_lines~5_combout ;
wire \data_num_lines~6_combout ;
wire \data_num_lines~9_combout ;
wire \data_num_lines~4_combout ;
wire \Selector18~4_combout ;
wire \Selector1~0_combout ;
wire \addr_num_lines~6_combout ;
wire \addr_num_lines~7_combout ;
wire \addr_num_lines~8_combout ;
wire \Equal0~0_combout ;
wire \addr_mem~0_combout ;
wire \addr_mem[1][0]~q ;
wire \addr_mem~1_combout ;
wire \addr_mem[2][0]~q ;
wire \addr_mem~2_combout ;
wire \addr_mem[0][0]~q ;
wire \Selector16~0_combout ;
wire \addr_mem~3_combout ;
wire \addr_mem[3][0]~q ;
wire \Selector16~1_combout ;
wire \header_information[0]~q ;
wire \Selector16~2_combout ;
wire \addr_mem~4_combout ;
wire \addr_mem[1][4]~q ;
wire \addr_mem~5_combout ;
wire \addr_mem[2][4]~q ;
wire \addr_mem~6_combout ;
wire \addr_mem[0][4]~q ;
wire \Selector12~0_combout ;
wire \addr_mem~7_combout ;
wire \addr_mem[3][4]~q ;
wire \Selector12~1_combout ;
wire \header_information[4]~q ;
wire \Selector12~2_combout ;
wire \addr_mem~8_combout ;
wire \addr_mem[1][2]~q ;
wire \addr_mem~9_combout ;
wire \addr_mem[2][2]~q ;
wire \addr_mem~10_combout ;
wire \addr_mem[0][2]~q ;
wire \Selector14~0_combout ;
wire \addr_mem~11_combout ;
wire \addr_mem[3][2]~q ;
wire \Selector14~1_combout ;
wire \header_information[2]~q ;
wire \Selector14~2_combout ;
wire \addr_mem~12_combout ;
wire \addr_mem[2][1]~q ;
wire \addr_mem~13_combout ;
wire \addr_mem[1][1]~q ;
wire \addr_mem~14_combout ;
wire \addr_mem[0][1]~q ;
wire \Selector15~0_combout ;
wire \addr_mem~15_combout ;
wire \addr_mem[3][1]~q ;
wire \Selector15~1_combout ;
wire \header_information[1]~q ;
wire \Selector9~0_combout ;
wire \Selector15~2_combout ;
wire \addr_mem~16_combout ;
wire \addr_mem[2][3]~q ;
wire \addr_mem~17_combout ;
wire \addr_mem[1][3]~q ;
wire \addr_mem~18_combout ;
wire \addr_mem[0][3]~q ;
wire \Selector13~0_combout ;
wire \addr_mem~19_combout ;
wire \addr_mem[3][3]~q ;
wire \Selector13~1_combout ;
wire \header_information[3]~q ;
wire \Selector13~2_combout ;
wire \addr_mem~20_combout ;
wire \addr_mem[2][5]~q ;
wire \addr_mem~21_combout ;
wire \addr_mem[1][5]~q ;
wire \addr_mem~22_combout ;
wire \addr_mem[0][5]~q ;
wire \Selector11~0_combout ;
wire \addr_mem~23_combout ;
wire \addr_mem[3][5]~q ;
wire \Selector11~1_combout ;
wire \header_information[5]~q ;
wire \Selector11~2_combout ;
wire \addr_mem~24_combout ;
wire \addr_mem[1][6]~q ;
wire \addr_mem~25_combout ;
wire \addr_mem[2][6]~q ;
wire \addr_mem~26_combout ;
wire \addr_mem[0][6]~q ;
wire \Selector10~0_combout ;
wire \addr_mem~27_combout ;
wire \addr_mem[3][6]~q ;
wire \Selector10~1_combout ;
wire \header_information[6]~q ;
wire \Selector10~2_combout ;
wire \addr_mem~28_combout ;
wire \addr_mem[2][7]~q ;
wire \addr_mem~29_combout ;
wire \addr_mem[1][7]~q ;
wire \addr_mem~30_combout ;
wire \addr_mem[0][7]~q ;
wire \Selector9~1_combout ;
wire \addr_mem~31_combout ;
wire \addr_mem[3][7]~q ;
wire \Selector9~2_combout ;
wire \header_information[7]~q ;
wire \Selector9~3_combout ;
wire \Selector3~5_combout ;


flashLoader_data_adapter_8_32 data_adapter_8_32_inst(
	.out_valid1(out_valid),
	.out_endofpacket1(out_endofpacket),
	.in_cmd_channel_reg_1(in_cmd_channel_reg_1),
	.stateST_WAIT_RSP(stateST_WAIT_RSP),
	.out_data_0(out_data_0),
	.out_data_1(\data_adapter_8_32_inst|out_data[1]~q ),
	.out_data_2(\data_adapter_8_32_inst|out_data[2]~q ),
	.out_data_3(\data_adapter_8_32_inst|out_data[3]~q ),
	.out_data_4(\data_adapter_8_32_inst|out_data[4]~q ),
	.out_data_5(\data_adapter_8_32_inst|out_data[5]~q ),
	.out_data_6(\data_adapter_8_32_inst|out_data[6]~q ),
	.out_data_7(\data_adapter_8_32_inst|out_data[7]~q ),
	.out_data_8(\data_adapter_8_32_inst|out_data[8]~q ),
	.out_data_9(\data_adapter_8_32_inst|out_data[9]~q ),
	.out_data_10(\data_adapter_8_32_inst|out_data[10]~q ),
	.out_data_11(\data_adapter_8_32_inst|out_data[11]~q ),
	.out_data_12(\data_adapter_8_32_inst|out_data[12]~q ),
	.out_data_13(\data_adapter_8_32_inst|out_data[13]~q ),
	.out_data_14(\data_adapter_8_32_inst|out_data[14]~q ),
	.out_data_15(\data_adapter_8_32_inst|out_data[15]~q ),
	.out_data_16(\data_adapter_8_32_inst|out_data[16]~q ),
	.out_data_17(\data_adapter_8_32_inst|out_data[17]~q ),
	.out_data_18(\data_adapter_8_32_inst|out_data[18]~q ),
	.out_data_19(\data_adapter_8_32_inst|out_data[19]~q ),
	.out_data_20(\data_adapter_8_32_inst|out_data[20]~q ),
	.out_data_21(\data_adapter_8_32_inst|out_data[21]~q ),
	.out_data_22(\data_adapter_8_32_inst|out_data[22]~q ),
	.out_data_23(\data_adapter_8_32_inst|out_data[23]~q ),
	.out_data_24(\data_adapter_8_32_inst|out_data[24]~q ),
	.out_data_25(\data_adapter_8_32_inst|out_data[25]~q ),
	.out_data_26(\data_adapter_8_32_inst|out_data[26]~q ),
	.out_data_27(\data_adapter_8_32_inst|out_data[27]~q ),
	.out_data_28(\data_adapter_8_32_inst|out_data[28]~q ),
	.out_data_29(\data_adapter_8_32_inst|out_data[29]~q ),
	.out_data_30(\data_adapter_8_32_inst|out_data[30]~q ),
	.out_data_31(\data_adapter_8_32_inst|out_data[31]~q ),
	.in_cmd_channel_reg_0(in_cmd_channel_reg_0),
	.a_valid1(\data_adapter_8_32_inst|a_valid~q ),
	.a_ready1(\data_adapter_8_32_inst|a_ready~combout ),
	.reset(\comb~0_combout ),
	.in_valid(\comb~1_combout ),
	.in_ready1(\data_adapter_8_32_inst|in_ready~combout ),
	.in_endofpacket(\in_rsp_eop~combout ),
	.in_data({out_rsp_data_71,out_rsp_data_61,out_rsp_data_51,out_rsp_data_41,out_rsp_data_32,out_rsp_data_210,out_rsp_data_110,out_rsp_data_01}),
	.clk(clk_clk));

flashLoader_data_adapter_32_8 data_adapter_32_8_inst(
	.reset(\comb~0_combout ),
	.state_register_1(\data_adapter_32_8_inst|state_register[1]~q ),
	.state_register_0(\data_adapter_32_8_inst|state_register[0]~q ),
	.out_valid1(\data_adapter_32_8_inst|out_valid~q ),
	.a_valid1(\data_adapter_32_8_inst|a_valid~q ),
	.stateST_SEND_DATA(stateST_SEND_DATA),
	.WideOr0(WideOr01),
	.WideOr01(WideOr04),
	.in_valid(\adap_in_cmd_valid~0_combout ),
	.out_data_0(\data_adapter_32_8_inst|out_data[0]~q ),
	.out_data_4(\data_adapter_32_8_inst|out_data[4]~q ),
	.out_data_2(\data_adapter_32_8_inst|out_data[2]~q ),
	.out_data_1(\data_adapter_32_8_inst|out_data[1]~q ),
	.out_data_3(\data_adapter_32_8_inst|out_data[3]~q ),
	.out_data_5(\data_adapter_32_8_inst|out_data[5]~q ),
	.out_data_6(\data_adapter_32_8_inst|out_data[6]~q ),
	.out_data_7(\data_adapter_32_8_inst|out_data[7]~q ),
	.in_data({\adap_in_cmd_data[31]~36_combout ,\adap_in_cmd_data[30]~29_combout ,\adap_in_cmd_data[29]~25_combout ,\adap_in_cmd_data[28]~9_combout ,\adap_in_cmd_data[27]~21_combout ,\adap_in_cmd_data[26]~13_combout ,\adap_in_cmd_data[25]~17_combout ,
\adap_in_cmd_data[24]~3_combout ,\adap_in_cmd_data[23]~30_combout ,\adap_in_cmd_data[22]~27_combout ,\adap_in_cmd_data[21]~22_combout ,\adap_in_cmd_data[20]~7_combout ,\adap_in_cmd_data[19]~18_combout ,\adap_in_cmd_data[18]~11_combout ,
\adap_in_cmd_data[17]~14_combout ,\adap_in_cmd_data[16]~1_combout ,\adap_in_cmd_data[15]~31_combout ,\adap_in_cmd_data[14]~26_combout ,\adap_in_cmd_data[13]~23_combout ,\adap_in_cmd_data[12]~6_combout ,\adap_in_cmd_data[11]~19_combout ,
\adap_in_cmd_data[10]~10_combout ,\adap_in_cmd_data[9]~15_combout ,\adap_in_cmd_data[8]~0_combout ,\adap_in_cmd_data[7]~32_combout ,\adap_in_cmd_data[6]~28_combout ,\adap_in_cmd_data[5]~24_combout ,\adap_in_cmd_data[4]~8_combout ,\adap_in_cmd_data[3]~20_combout ,
\adap_in_cmd_data[2]~12_combout ,\adap_in_cmd_data[1]~16_combout ,\adap_in_cmd_data[0]~2_combout }),
	.clk(clk_clk));

cycloneive_lcell_comb \comb~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(reset),
	.datad(stateST_IDLE),
	.cin(gnd),
	.combout(\comb~0_combout ),
	.cout());
defparam \comb~0 .lut_mask = 16'h0FFF;
defparam \comb~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \comb~1 (
	.dataa(out_rsp_valid),
	.datab(\state.ST_WAIT_RSP~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\comb~1_combout ),
	.cout());
defparam \comb~1 .lut_mask = 16'h8888;
defparam \comb~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_valid~0 (
	.dataa(WideOr1),
	.datab(stateST_SEND_DATA),
	.datac(stateST_SEND_ADDR),
	.datad(gnd),
	.cin(gnd),
	.combout(\adap_in_cmd_valid~0_combout ),
	.cout());
defparam \adap_in_cmd_valid~0 .lut_mask = 16'hA8A8;
defparam \adap_in_cmd_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[8]~0 (
	.dataa(src_data_8),
	.datab(in_cmd_channel[0]),
	.datac(cmd_data_8),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[8]~0_combout ),
	.cout());
defparam \adap_in_cmd_data[8]~0 .lut_mask = 16'h00EA;
defparam \adap_in_cmd_data[8]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[16]~1 (
	.dataa(src_data_16),
	.datab(in_cmd_channel[0]),
	.datac(src_data_161),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[16]~1_combout ),
	.cout());
defparam \adap_in_cmd_data[16]~1 .lut_mask = 16'h00EA;
defparam \adap_in_cmd_data[16]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[0]~2 (
	.dataa(in_cmd_data[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[0]~2_combout ),
	.cout());
defparam \adap_in_cmd_data[0]~2 .lut_mask = 16'h00AA;
defparam \adap_in_cmd_data[0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[24]~3 (
	.dataa(in_cmd_data[24]),
	.datab(gnd),
	.datac(gnd),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[24]~3_combout ),
	.cout());
defparam \adap_in_cmd_data[24]~3 .lut_mask = 16'h00AA;
defparam \adap_in_cmd_data[24]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[12]~4 (
	.dataa(csr_flash_cmd_wr_data_0_data_12),
	.datab(stateST_SEND_HEADER),
	.datac(has_dummy),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\adap_in_cmd_data[12]~4_combout ),
	.cout());
defparam \adap_in_cmd_data[12]~4 .lut_mask = 16'hAAC0;
defparam \adap_in_cmd_data[12]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[12]~5 (
	.dataa(in_cmd_channel[1]),
	.datab(csr_flash_cmd_wr_data_1_data_12),
	.datac(\adap_in_cmd_data[12]~4_combout ),
	.datad(stateST_SEND_DATA_1),
	.cin(gnd),
	.combout(\adap_in_cmd_data[12]~5_combout ),
	.cout());
defparam \adap_in_cmd_data[12]~5 .lut_mask = 16'h88A0;
defparam \adap_in_cmd_data[12]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[12]~6 (
	.dataa(\adap_in_cmd_data[12]~5_combout ),
	.datab(in_cmd_channel[0]),
	.datac(cmd_data_12),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[12]~6_combout ),
	.cout());
defparam \adap_in_cmd_data[12]~6 .lut_mask = 16'h00EA;
defparam \adap_in_cmd_data[12]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[20]~7 (
	.dataa(src_data_20),
	.datab(in_cmd_channel[0]),
	.datac(src_data_201),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[20]~7_combout ),
	.cout());
defparam \adap_in_cmd_data[20]~7 .lut_mask = 16'h00EA;
defparam \adap_in_cmd_data[20]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[4]~8 (
	.dataa(in_cmd_data[4]),
	.datab(gnd),
	.datac(gnd),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[4]~8_combout ),
	.cout());
defparam \adap_in_cmd_data[4]~8 .lut_mask = 16'h00AA;
defparam \adap_in_cmd_data[4]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[28]~9 (
	.dataa(src_data_28),
	.datab(in_cmd_channel[0]),
	.datac(src_data_281),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[28]~9_combout ),
	.cout());
defparam \adap_in_cmd_data[28]~9 .lut_mask = 16'h00EA;
defparam \adap_in_cmd_data[28]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[10]~10 (
	.dataa(src_data_10),
	.datab(in_cmd_channel[0]),
	.datac(cmd_data_10),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[10]~10_combout ),
	.cout());
defparam \adap_in_cmd_data[10]~10 .lut_mask = 16'h00EA;
defparam \adap_in_cmd_data[10]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[18]~11 (
	.dataa(in_cmd_data[18]),
	.datab(gnd),
	.datac(gnd),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[18]~11_combout ),
	.cout());
defparam \adap_in_cmd_data[18]~11 .lut_mask = 16'h00AA;
defparam \adap_in_cmd_data[18]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[2]~12 (
	.dataa(in_cmd_data[2]),
	.datab(gnd),
	.datac(gnd),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[2]~12_combout ),
	.cout());
defparam \adap_in_cmd_data[2]~12 .lut_mask = 16'h00AA;
defparam \adap_in_cmd_data[2]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[26]~13 (
	.dataa(in_cmd_data[26]),
	.datab(gnd),
	.datac(gnd),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[26]~13_combout ),
	.cout());
defparam \adap_in_cmd_data[26]~13 .lut_mask = 16'h00AA;
defparam \adap_in_cmd_data[26]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[17]~14 (
	.dataa(src_data_17),
	.datab(in_cmd_channel[0]),
	.datac(src_data_171),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[17]~14_combout ),
	.cout());
defparam \adap_in_cmd_data[17]~14 .lut_mask = 16'h00EA;
defparam \adap_in_cmd_data[17]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[9]~15 (
	.dataa(src_data_9),
	.datab(in_cmd_channel[0]),
	.datac(cmd_data_9),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[9]~15_combout ),
	.cout());
defparam \adap_in_cmd_data[9]~15 .lut_mask = 16'h00EA;
defparam \adap_in_cmd_data[9]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[1]~16 (
	.dataa(in_cmd_data[1]),
	.datab(gnd),
	.datac(gnd),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[1]~16_combout ),
	.cout());
defparam \adap_in_cmd_data[1]~16 .lut_mask = 16'h00AA;
defparam \adap_in_cmd_data[1]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[25]~17 (
	.dataa(in_cmd_data[25]),
	.datab(gnd),
	.datac(gnd),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[25]~17_combout ),
	.cout());
defparam \adap_in_cmd_data[25]~17 .lut_mask = 16'h00AA;
defparam \adap_in_cmd_data[25]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[19]~18 (
	.dataa(src_data_19),
	.datab(src_data_191),
	.datac(gnd),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[19]~18_combout ),
	.cout());
defparam \adap_in_cmd_data[19]~18 .lut_mask = 16'h00EE;
defparam \adap_in_cmd_data[19]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[11]~19 (
	.dataa(src_data_11),
	.datab(in_cmd_channel[0]),
	.datac(cmd_data_11),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[11]~19_combout ),
	.cout());
defparam \adap_in_cmd_data[11]~19 .lut_mask = 16'h00EA;
defparam \adap_in_cmd_data[11]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[3]~20 (
	.dataa(in_cmd_data[3]),
	.datab(gnd),
	.datac(gnd),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[3]~20_combout ),
	.cout());
defparam \adap_in_cmd_data[3]~20 .lut_mask = 16'h00AA;
defparam \adap_in_cmd_data[3]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[27]~21 (
	.dataa(src_data_27),
	.datab(in_cmd_channel[0]),
	.datac(src_data_271),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[27]~21_combout ),
	.cout());
defparam \adap_in_cmd_data[27]~21 .lut_mask = 16'h00EA;
defparam \adap_in_cmd_data[27]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[21]~22 (
	.dataa(src_data_21),
	.datab(in_cmd_channel[0]),
	.datac(src_data_211),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[21]~22_combout ),
	.cout());
defparam \adap_in_cmd_data[21]~22 .lut_mask = 16'h00EA;
defparam \adap_in_cmd_data[21]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[13]~23 (
	.dataa(src_data_13),
	.datab(in_cmd_channel[0]),
	.datac(cmd_data_13),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[13]~23_combout ),
	.cout());
defparam \adap_in_cmd_data[13]~23 .lut_mask = 16'h00EA;
defparam \adap_in_cmd_data[13]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[5]~24 (
	.dataa(in_cmd_data[5]),
	.datab(gnd),
	.datac(gnd),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[5]~24_combout ),
	.cout());
defparam \adap_in_cmd_data[5]~24 .lut_mask = 16'h00AA;
defparam \adap_in_cmd_data[5]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[29]~25 (
	.dataa(src_data_29),
	.datab(in_cmd_channel[0]),
	.datac(src_data_291),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[29]~25_combout ),
	.cout());
defparam \adap_in_cmd_data[29]~25 .lut_mask = 16'h00EA;
defparam \adap_in_cmd_data[29]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[14]~26 (
	.dataa(src_data_14),
	.datab(in_cmd_channel[0]),
	.datac(cmd_data_14),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[14]~26_combout ),
	.cout());
defparam \adap_in_cmd_data[14]~26 .lut_mask = 16'h00EA;
defparam \adap_in_cmd_data[14]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[22]~27 (
	.dataa(in_cmd_data[22]),
	.datab(gnd),
	.datac(gnd),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[22]~27_combout ),
	.cout());
defparam \adap_in_cmd_data[22]~27 .lut_mask = 16'h00AA;
defparam \adap_in_cmd_data[22]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[6]~28 (
	.dataa(in_cmd_data[6]),
	.datab(gnd),
	.datac(gnd),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[6]~28_combout ),
	.cout());
defparam \adap_in_cmd_data[6]~28 .lut_mask = 16'h00AA;
defparam \adap_in_cmd_data[6]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[30]~29 (
	.dataa(src_data_30),
	.datab(in_cmd_channel[0]),
	.datac(src_data_302),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[30]~29_combout ),
	.cout());
defparam \adap_in_cmd_data[30]~29 .lut_mask = 16'h00EA;
defparam \adap_in_cmd_data[30]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[23]~30 (
	.dataa(in_cmd_data[23]),
	.datab(gnd),
	.datac(gnd),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[23]~30_combout ),
	.cout());
defparam \adap_in_cmd_data[23]~30 .lut_mask = 16'h00AA;
defparam \adap_in_cmd_data[23]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[15]~31 (
	.dataa(src_data_15),
	.datab(in_cmd_channel[0]),
	.datac(cmd_data_15),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[15]~31_combout ),
	.cout());
defparam \adap_in_cmd_data[15]~31 .lut_mask = 16'h00EA;
defparam \adap_in_cmd_data[15]~31 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[7]~32 (
	.dataa(in_cmd_data[7]),
	.datab(gnd),
	.datac(gnd),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[7]~32_combout ),
	.cout());
defparam \adap_in_cmd_data[7]~32 .lut_mask = 16'h00AA;
defparam \adap_in_cmd_data[7]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[31]~33 (
	.dataa(is_burst_reg),
	.datab(src_data_301),
	.datac(mem_write_data_reg_31),
	.datad(out_payload_31),
	.cin(gnd),
	.combout(\adap_in_cmd_data[31]~33_combout ),
	.cout());
defparam \adap_in_cmd_data[31]~33 .lut_mask = 16'hEAC0;
defparam \adap_in_cmd_data[31]~33 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[31]~34 (
	.dataa(in_cmd_channel[0]),
	.datab(current_stateSTATE_WR_DATA),
	.datac(\adap_in_cmd_data[31]~33_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\adap_in_cmd_data[31]~34_combout ),
	.cout());
defparam \adap_in_cmd_data[31]~34 .lut_mask = 16'h8080;
defparam \adap_in_cmd_data[31]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[31]~35 (
	.dataa(csr_flash_cmd_wr_data_0_data_31),
	.datab(csr_flash_cmd_wr_data_1_data_31),
	.datac(stateST_SEND_DATA_1),
	.datad(stateST_SEND_DATA_0),
	.cin(gnd),
	.combout(\adap_in_cmd_data[31]~35_combout ),
	.cout());
defparam \adap_in_cmd_data[31]~35 .lut_mask = 16'hEAC0;
defparam \adap_in_cmd_data[31]~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \adap_in_cmd_data[31]~36 (
	.dataa(\adap_in_cmd_data[31]~34_combout ),
	.datab(in_cmd_channel[1]),
	.datac(\adap_in_cmd_data[31]~35_combout ),
	.datad(src_startofpacket),
	.cin(gnd),
	.combout(\adap_in_cmd_data[31]~36_combout ),
	.cout());
defparam \adap_in_cmd_data[31]~36 .lut_mask = 16'h00EA;
defparam \adap_in_cmd_data[31]~36 .sum_lutc_input = "datac";

dffeas \data_num_lines[1] (
	.clk(clk_clk),
	.d(\data_num_lines[1]~0_combout ),
	.asdata(\Equal3~0_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always2~1_combout ),
	.ena(\always0~1_combout ),
	.q(data_num_lines_1),
	.prn(vcc));
defparam \data_num_lines[1] .is_wysiwyg = "true";
defparam \data_num_lines[1] .power_up = "low";

dffeas \data_num_lines[2] (
	.clk(clk_clk),
	.d(\data_num_lines[2]~1_combout ),
	.asdata(\Equal4~0_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always2~1_combout ),
	.ena(\always0~1_combout ),
	.q(data_num_lines_2),
	.prn(vcc));
defparam \data_num_lines[2] .is_wysiwyg = "true";
defparam \data_num_lines[2] .power_up = "low";

dffeas \addr_num_lines[2] (
	.clk(clk_clk),
	.d(\addr_num_lines[2]~1_combout ),
	.asdata(\Equal4~0_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always2~1_combout ),
	.ena(\always0~1_combout ),
	.q(addr_num_lines_2),
	.prn(vcc));
defparam \addr_num_lines[2] .is_wysiwyg = "true";
defparam \addr_num_lines[2] .power_up = "low";

dffeas \addr_num_lines[1] (
	.clk(clk_clk),
	.d(\addr_num_lines[1]~0_combout ),
	.asdata(\Equal3~0_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always2~1_combout ),
	.ena(\always0~1_combout ),
	.q(addr_num_lines_1),
	.prn(vcc));
defparam \addr_num_lines[1] .is_wysiwyg = "true";
defparam \addr_num_lines[1] .power_up = "low";

dffeas \state.ST_SEND_DUMMY_RSP (
	.clk(clk_clk),
	.d(\Selector6~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stateST_SEND_DUMMY_RSP),
	.prn(vcc));
defparam \state.ST_SEND_DUMMY_RSP .is_wysiwyg = "true";
defparam \state.ST_SEND_DUMMY_RSP .power_up = "low";

dffeas \in_cmd_channel_reg[1] (
	.clk(clk_clk),
	.d(in_cmd_channel[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(in_cmd_channel_reg_1),
	.prn(vcc));
defparam \in_cmd_channel_reg[1] .is_wysiwyg = "true";
defparam \in_cmd_channel_reg[1] .power_up = "low";

cycloneive_lcell_comb \out_rsp_data[0]~0 (
	.dataa(out_valid),
	.datab(out_data_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_0),
	.cout());
defparam \out_rsp_data[0]~0 .lut_mask = 16'h8888;
defparam \out_rsp_data[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[1]~1 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_1),
	.cout());
defparam \out_rsp_data[1]~1 .lut_mask = 16'h8888;
defparam \out_rsp_data[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[2]~2 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_2),
	.cout());
defparam \out_rsp_data[2]~2 .lut_mask = 16'h8888;
defparam \out_rsp_data[2]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[3]~3 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_3),
	.cout());
defparam \out_rsp_data[3]~3 .lut_mask = 16'h8888;
defparam \out_rsp_data[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[4]~4 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_4),
	.cout());
defparam \out_rsp_data[4]~4 .lut_mask = 16'h8888;
defparam \out_rsp_data[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[5]~5 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_5),
	.cout());
defparam \out_rsp_data[5]~5 .lut_mask = 16'h8888;
defparam \out_rsp_data[5]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[6]~6 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_6),
	.cout());
defparam \out_rsp_data[6]~6 .lut_mask = 16'h8888;
defparam \out_rsp_data[6]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[7]~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(out_valid),
	.datad(\data_adapter_8_32_inst|out_data[7]~q ),
	.cin(gnd),
	.combout(out_rsp_data_7),
	.cout());
defparam \out_rsp_data[7]~7 .lut_mask = 16'hF000;
defparam \out_rsp_data[7]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[8]~8 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_8),
	.cout());
defparam \out_rsp_data[8]~8 .lut_mask = 16'h8888;
defparam \out_rsp_data[8]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[9]~9 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_9),
	.cout());
defparam \out_rsp_data[9]~9 .lut_mask = 16'h8888;
defparam \out_rsp_data[9]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[10]~10 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_10),
	.cout());
defparam \out_rsp_data[10]~10 .lut_mask = 16'h8888;
defparam \out_rsp_data[10]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[11]~11 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_11),
	.cout());
defparam \out_rsp_data[11]~11 .lut_mask = 16'h8888;
defparam \out_rsp_data[11]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[12]~12 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_12),
	.cout());
defparam \out_rsp_data[12]~12 .lut_mask = 16'h8888;
defparam \out_rsp_data[12]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[13]~13 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_13),
	.cout());
defparam \out_rsp_data[13]~13 .lut_mask = 16'h8888;
defparam \out_rsp_data[13]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[14]~14 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_14),
	.cout());
defparam \out_rsp_data[14]~14 .lut_mask = 16'h8888;
defparam \out_rsp_data[14]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[15]~15 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_15),
	.cout());
defparam \out_rsp_data[15]~15 .lut_mask = 16'h8888;
defparam \out_rsp_data[15]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[16]~16 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[16]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_16),
	.cout());
defparam \out_rsp_data[16]~16 .lut_mask = 16'h8888;
defparam \out_rsp_data[16]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[17]~17 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[17]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_17),
	.cout());
defparam \out_rsp_data[17]~17 .lut_mask = 16'h8888;
defparam \out_rsp_data[17]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[18]~18 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[18]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_18),
	.cout());
defparam \out_rsp_data[18]~18 .lut_mask = 16'h8888;
defparam \out_rsp_data[18]~18 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[19]~19 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[19]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_19),
	.cout());
defparam \out_rsp_data[19]~19 .lut_mask = 16'h8888;
defparam \out_rsp_data[19]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[20]~20 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[20]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_20),
	.cout());
defparam \out_rsp_data[20]~20 .lut_mask = 16'h8888;
defparam \out_rsp_data[20]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[21]~21 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[21]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_21),
	.cout());
defparam \out_rsp_data[21]~21 .lut_mask = 16'h8888;
defparam \out_rsp_data[21]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[22]~22 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[22]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_22),
	.cout());
defparam \out_rsp_data[22]~22 .lut_mask = 16'h8888;
defparam \out_rsp_data[22]~22 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[23]~23 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[23]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_23),
	.cout());
defparam \out_rsp_data[23]~23 .lut_mask = 16'h8888;
defparam \out_rsp_data[23]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[24]~24 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[24]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_24),
	.cout());
defparam \out_rsp_data[24]~24 .lut_mask = 16'h8888;
defparam \out_rsp_data[24]~24 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[25]~25 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[25]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_25),
	.cout());
defparam \out_rsp_data[25]~25 .lut_mask = 16'h8888;
defparam \out_rsp_data[25]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[26]~26 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[26]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_26),
	.cout());
defparam \out_rsp_data[26]~26 .lut_mask = 16'h8888;
defparam \out_rsp_data[26]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[27]~27 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[27]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_27),
	.cout());
defparam \out_rsp_data[27]~27 .lut_mask = 16'h8888;
defparam \out_rsp_data[27]~27 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[28]~28 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[28]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_28),
	.cout());
defparam \out_rsp_data[28]~28 .lut_mask = 16'h8888;
defparam \out_rsp_data[28]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[29]~29 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[29]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_29),
	.cout());
defparam \out_rsp_data[29]~29 .lut_mask = 16'h8888;
defparam \out_rsp_data[29]~29 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[30]~30 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[30]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_30),
	.cout());
defparam \out_rsp_data[30]~30 .lut_mask = 16'h8888;
defparam \out_rsp_data[30]~30 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_rsp_data[31]~31 (
	.dataa(out_valid),
	.datab(\data_adapter_8_32_inst|out_data[31]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_rsp_data_31),
	.cout());
defparam \out_rsp_data[31]~31 .lut_mask = 16'h8888;
defparam \out_rsp_data[31]~31 .sum_lutc_input = "datac";

dffeas \in_cmd_channel_reg[0] (
	.clk(clk_clk),
	.d(in_cmd_channel[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(in_cmd_channel_reg_0),
	.prn(vcc));
defparam \in_cmd_channel_reg[0] .is_wysiwyg = "true";
defparam \in_cmd_channel_reg[0] .power_up = "low";

dffeas \header_information[30] (
	.clk(clk_clk),
	.d(in_cmd_data[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(header_information_30),
	.prn(vcc));
defparam \header_information[30] .is_wysiwyg = "true";
defparam \header_information[30] .power_up = "low";

dffeas \header_information[29] (
	.clk(clk_clk),
	.d(in_cmd_data[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(header_information_29),
	.prn(vcc));
defparam \header_information[29] .is_wysiwyg = "true";
defparam \header_information[29] .power_up = "low";

dffeas \header_information[28] (
	.clk(clk_clk),
	.d(in_cmd_data[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(header_information_28),
	.prn(vcc));
defparam \header_information[28] .is_wysiwyg = "true";
defparam \header_information[28] .power_up = "low";

dffeas \header_information[27] (
	.clk(clk_clk),
	.d(in_cmd_data[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(header_information_27),
	.prn(vcc));
defparam \header_information[27] .is_wysiwyg = "true";
defparam \header_information[27] .power_up = "low";

dffeas \state.ST_IDLE (
	.clk(clk_clk),
	.d(\Selector0~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stateST_IDLE),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

dffeas \state.ST_SEND_DATA (
	.clk(clk_clk),
	.d(\Selector3~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stateST_SEND_DATA),
	.prn(vcc));
defparam \state.ST_SEND_DATA .is_wysiwyg = "true";
defparam \state.ST_SEND_DATA .power_up = "low";

dffeas \state.ST_SEND_ADDR (
	.clk(clk_clk),
	.d(\Selector2~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stateST_SEND_ADDR),
	.prn(vcc));
defparam \state.ST_SEND_ADDR .is_wysiwyg = "true";
defparam \state.ST_SEND_ADDR .power_up = "low";

cycloneive_lcell_comb \Selector18~2 (
	.dataa(\Selector18~0_combout ),
	.datab(\Selector18~1_combout ),
	.datac(gnd),
	.datad(stateST_IDLE),
	.cin(gnd),
	.combout(Selector18),
	.cout());
defparam \Selector18~2 .lut_mask = 16'h88FF;
defparam \Selector18~2 .sum_lutc_input = "datac";

dffeas \op_num_lines[1] (
	.clk(clk_clk),
	.d(\Equal3~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(op_num_lines_1),
	.prn(vcc));
defparam \op_num_lines[1] .is_wysiwyg = "true";
defparam \op_num_lines[1] .power_up = "low";

dffeas \data_num_lines[0] (
	.clk(clk_clk),
	.d(\data_num_lines~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_num_lines_0),
	.prn(vcc));
defparam \data_num_lines[0] .is_wysiwyg = "true";
defparam \data_num_lines[0] .power_up = "low";

dffeas \op_num_lines[0] (
	.clk(clk_clk),
	.d(\data_num_lines~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(op_num_lines_0),
	.prn(vcc));
defparam \op_num_lines[0] .is_wysiwyg = "true";
defparam \op_num_lines[0] .power_up = "low";

dffeas \op_num_lines[2] (
	.clk(clk_clk),
	.d(\Equal4~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(op_num_lines_2),
	.prn(vcc));
defparam \op_num_lines[2] .is_wysiwyg = "true";
defparam \op_num_lines[2] .power_up = "low";

cycloneive_lcell_comb \adap_out_cmd_ready~0 (
	.dataa(stateST_SEND_DATA),
	.datab(WideOr01),
	.datac(in_ready),
	.datad(WideOr02),
	.cin(gnd),
	.combout(adap_out_cmd_ready),
	.cout());
defparam \adap_out_cmd_ready~0 .lut_mask = 16'hA888;
defparam \adap_out_cmd_ready~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector18~3 (
	.dataa(\data_adapter_32_8_inst|state_register[1]~q ),
	.datab(\data_adapter_32_8_inst|state_register[0]~q ),
	.datac(gnd),
	.datad(\last_word_detect~q ),
	.cin(gnd),
	.combout(Selector181),
	.cout());
defparam \Selector18~3 .lut_mask = 16'h0088;
defparam \Selector18~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector18~5 (
	.dataa(Selector181),
	.datab(stateST_SEND_DATA),
	.datac(Selector18),
	.datad(\Selector18~4_combout ),
	.cin(gnd),
	.combout(Selector182),
	.cout());
defparam \Selector18~5 .lut_mask = 16'hF8F0;
defparam \Selector18~5 .sum_lutc_input = "datac";

dffeas \header_information[11] (
	.clk(clk_clk),
	.d(in_cmd_data[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(header_information_11),
	.prn(vcc));
defparam \header_information[11] .is_wysiwyg = "true";
defparam \header_information[11] .power_up = "low";

dffeas \state.ST_SEND_OPCODE (
	.clk(clk_clk),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stateST_SEND_OPCODE),
	.prn(vcc));
defparam \state.ST_SEND_OPCODE .is_wysiwyg = "true";
defparam \state.ST_SEND_OPCODE .power_up = "low";

cycloneive_lcell_comb \Selector8~0 (
	.dataa(stateST_SEND_ADDR),
	.datab(stateST_SEND_OPCODE),
	.datac(stateST_SEND_DATA),
	.datad(\data_adapter_32_8_inst|out_valid~q ),
	.cin(gnd),
	.combout(Selector8),
	.cout());
defparam \Selector8~0 .lut_mask = 16'hFEEE;
defparam \Selector8~0 .sum_lutc_input = "datac";

dffeas \addr_num_lines[0] (
	.clk(clk_clk),
	.d(\addr_num_lines~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(addr_num_lines_0),
	.prn(vcc));
defparam \addr_num_lines[0] .is_wysiwyg = "true";
defparam \addr_num_lines[0] .power_up = "low";

dffeas \header_information[13] (
	.clk(clk_clk),
	.d(in_cmd_data[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(header_information_13),
	.prn(vcc));
defparam \header_information[13] .is_wysiwyg = "true";
defparam \header_information[13] .power_up = "low";

dffeas \header_information[17] (
	.clk(clk_clk),
	.d(in_cmd_data[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(header_information_17),
	.prn(vcc));
defparam \header_information[17] .is_wysiwyg = "true";
defparam \header_information[17] .power_up = "low";

dffeas \header_information[16] (
	.clk(clk_clk),
	.d(in_cmd_data[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(header_information_16),
	.prn(vcc));
defparam \header_information[16] .is_wysiwyg = "true";
defparam \header_information[16] .power_up = "low";

dffeas \header_information[15] (
	.clk(clk_clk),
	.d(in_cmd_data[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(header_information_15),
	.prn(vcc));
defparam \header_information[15] .is_wysiwyg = "true";
defparam \header_information[15] .power_up = "low";

dffeas \header_information[14] (
	.clk(clk_clk),
	.d(in_cmd_data[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(header_information_14),
	.prn(vcc));
defparam \header_information[14] .is_wysiwyg = "true";
defparam \header_information[14] .power_up = "low";

cycloneive_lcell_comb \Selector20~2 (
	.dataa(stateST_SEND_OPCODE),
	.datab(\Selector20~1_combout ),
	.datac(stateST_SEND_DATA),
	.datad(\data_in_cnt_done~combout ),
	.cin(gnd),
	.combout(Selector20),
	.cout());
defparam \Selector20~2 .lut_mask = 16'hFEEE;
defparam \Selector20~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector16~3 (
	.dataa(\data_adapter_32_8_inst|out_data[0]~q ),
	.datab(\Selector16~2_combout ),
	.datac(gnd),
	.datad(stateST_SEND_DATA),
	.cin(gnd),
	.combout(Selector16),
	.cout());
defparam \Selector16~3 .lut_mask = 16'hAACC;
defparam \Selector16~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector12~3 (
	.dataa(\data_adapter_32_8_inst|out_data[4]~q ),
	.datab(\Selector12~2_combout ),
	.datac(gnd),
	.datad(stateST_SEND_DATA),
	.cin(gnd),
	.combout(Selector12),
	.cout());
defparam \Selector12~3 .lut_mask = 16'hAACC;
defparam \Selector12~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector14~3 (
	.dataa(\data_adapter_32_8_inst|out_data[2]~q ),
	.datab(\Selector14~2_combout ),
	.datac(gnd),
	.datad(stateST_SEND_DATA),
	.cin(gnd),
	.combout(Selector14),
	.cout());
defparam \Selector14~3 .lut_mask = 16'hAACC;
defparam \Selector14~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector15~3 (
	.dataa(\Selector15~2_combout ),
	.datab(stateST_SEND_DATA),
	.datac(\data_adapter_32_8_inst|out_data[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(Selector15),
	.cout());
defparam \Selector15~3 .lut_mask = 16'hEAEA;
defparam \Selector15~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector13~3 (
	.dataa(\Selector13~2_combout ),
	.datab(stateST_SEND_DATA),
	.datac(\data_adapter_32_8_inst|out_data[3]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(Selector13),
	.cout());
defparam \Selector13~3 .lut_mask = 16'hEAEA;
defparam \Selector13~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector11~3 (
	.dataa(\Selector11~2_combout ),
	.datab(stateST_SEND_DATA),
	.datac(\data_adapter_32_8_inst|out_data[5]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(Selector11),
	.cout());
defparam \Selector11~3 .lut_mask = 16'hEAEA;
defparam \Selector11~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector10~3 (
	.dataa(\data_adapter_32_8_inst|out_data[6]~q ),
	.datab(\Selector10~2_combout ),
	.datac(gnd),
	.datad(stateST_SEND_DATA),
	.cin(gnd),
	.combout(Selector10),
	.cout());
defparam \Selector10~3 .lut_mask = 16'hAACC;
defparam \Selector10~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector9~4 (
	.dataa(\Selector9~3_combout ),
	.datab(stateST_SEND_DATA),
	.datac(\data_adapter_32_8_inst|out_data[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(Selector9),
	.cout());
defparam \Selector9~4 .lut_mask = 16'hEAEA;
defparam \Selector9~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector17~0 (
	.dataa(\Selector4~0_combout ),
	.datab(\Selector3~5_combout ),
	.datac(\Selector20~1_combout ),
	.datad(\header_information[10]~q ),
	.cin(gnd),
	.combout(Selector17),
	.cout());
defparam \Selector17~0 .lut_mask = 16'hAAFE;
defparam \Selector17~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal12~0 (
	.dataa(csr_op_protocol_data_16),
	.datab(gnd),
	.datac(gnd),
	.datad(csr_op_protocol_data_17),
	.cin(gnd),
	.combout(\Equal12~0_combout ),
	.cout());
defparam \Equal12~0 .lut_mask = 16'h00AA;
defparam \Equal12~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal8~0 (
	.dataa(csr_op_protocol_data_8),
	.datab(gnd),
	.datac(gnd),
	.datad(csr_op_protocol_data_9),
	.cin(gnd),
	.combout(\Equal8~0_combout ),
	.cout());
defparam \Equal8~0 .lut_mask = 16'h00AA;
defparam \Equal8~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal5~0 (
	.dataa(current_stateSTATE_WR_DATA),
	.datab(current_stateSTATE_WR_CMD),
	.datac(current_stateSTATE_READ_DATA),
	.datad(current_stateSTATE_READ_CMD),
	.cin(gnd),
	.combout(\Equal5~0_combout ),
	.cout());
defparam \Equal5~0 .lut_mask = 16'h000E;
defparam \Equal5~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_num_lines[1]~0 (
	.dataa(\Equal12~0_combout ),
	.datab(\Equal8~0_combout ),
	.datac(gnd),
	.datad(\Equal5~0_combout ),
	.cin(gnd),
	.combout(\data_num_lines[1]~0_combout ),
	.cout());
defparam \data_num_lines[1]~0 .lut_mask = 16'hCCAA;
defparam \data_num_lines[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal3~0 (
	.dataa(csr_op_protocol_data_0),
	.datab(gnd),
	.datac(gnd),
	.datad(csr_op_protocol_data_1),
	.cin(gnd),
	.combout(\Equal3~0_combout ),
	.cout());
defparam \Equal3~0 .lut_mask = 16'h00AA;
defparam \Equal3~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always2~0 (
	.dataa(current_stateSTATE_READ_DATA),
	.datab(current_stateSTATE_WR_DATA),
	.datac(current_stateSTATE_WR_CMD),
	.datad(current_stateSTATE_READ_CMD),
	.cin(gnd),
	.combout(\always2~0_combout ),
	.cout());
defparam \always2~0 .lut_mask = 16'h0001;
defparam \always2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always2~1 (
	.dataa(\always2~0_combout ),
	.datab(gnd),
	.datac(in_cmd_channel[1]),
	.datad(in_cmd_channel[0]),
	.cin(gnd),
	.combout(\always2~1_combout ),
	.cout());
defparam \always2~1 .lut_mask = 16'h0AF0;
defparam \always2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always0~0 (
	.dataa(src_startofpacket),
	.datab(src_valid),
	.datac(in_cmd_channel[0]),
	.datad(cmd_valid),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
defparam \always0~0 .lut_mask = 16'hA888;
defparam \always0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always0~1 (
	.dataa(\always0~0_combout ),
	.datab(Selector18),
	.datac(adap_out_cmd_ready),
	.datad(Selector181),
	.cin(gnd),
	.combout(\always0~1_combout ),
	.cout());
defparam \always0~1 .lut_mask = 16'hA888;
defparam \always0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_num_lines~7 (
	.dataa(csr_op_protocol_data_17),
	.datab(gnd),
	.datac(gnd),
	.datad(csr_op_protocol_data_16),
	.cin(gnd),
	.combout(\data_num_lines~7_combout ),
	.cout());
defparam \data_num_lines~7 .lut_mask = 16'h00AA;
defparam \data_num_lines~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_num_lines~8 (
	.dataa(csr_op_protocol_data_9),
	.datab(gnd),
	.datac(gnd),
	.datad(csr_op_protocol_data_8),
	.cin(gnd),
	.combout(\data_num_lines~8_combout ),
	.cout());
defparam \data_num_lines~8 .lut_mask = 16'h00AA;
defparam \data_num_lines~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_num_lines[2]~1 (
	.dataa(\data_num_lines~7_combout ),
	.datab(\data_num_lines~8_combout ),
	.datac(gnd),
	.datad(\Equal5~0_combout ),
	.cin(gnd),
	.combout(\data_num_lines[2]~1_combout ),
	.cout());
defparam \data_num_lines[2]~1 .lut_mask = 16'hCCAA;
defparam \data_num_lines[2]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal4~0 (
	.dataa(csr_op_protocol_data_1),
	.datab(gnd),
	.datac(gnd),
	.datad(csr_op_protocol_data_0),
	.cin(gnd),
	.combout(\Equal4~0_combout ),
	.cout());
defparam \Equal4~0 .lut_mask = 16'h00AA;
defparam \Equal4~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_num_lines~4 (
	.dataa(csr_op_protocol_data_13),
	.datab(gnd),
	.datac(gnd),
	.datad(csr_op_protocol_data_12),
	.cin(gnd),
	.combout(\addr_num_lines~4_combout ),
	.cout());
defparam \addr_num_lines~4 .lut_mask = 16'h00AA;
defparam \addr_num_lines~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_num_lines~5 (
	.dataa(csr_op_protocol_data_5),
	.datab(gnd),
	.datac(gnd),
	.datad(csr_op_protocol_data_4),
	.cin(gnd),
	.combout(\addr_num_lines~5_combout ),
	.cout());
defparam \addr_num_lines~5 .lut_mask = 16'h00AA;
defparam \addr_num_lines~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_num_lines[2]~1 (
	.dataa(\addr_num_lines~4_combout ),
	.datab(\addr_num_lines~5_combout ),
	.datac(gnd),
	.datad(\Equal5~0_combout ),
	.cin(gnd),
	.combout(\addr_num_lines[2]~1_combout ),
	.cout());
defparam \addr_num_lines[2]~1 .lut_mask = 16'hCCAA;
defparam \addr_num_lines[2]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal10~0 (
	.dataa(csr_op_protocol_data_12),
	.datab(gnd),
	.datac(gnd),
	.datad(csr_op_protocol_data_13),
	.cin(gnd),
	.combout(\Equal10~0_combout ),
	.cout());
defparam \Equal10~0 .lut_mask = 16'h00AA;
defparam \Equal10~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal6~0 (
	.dataa(csr_op_protocol_data_4),
	.datab(gnd),
	.datac(gnd),
	.datad(csr_op_protocol_data_5),
	.cin(gnd),
	.combout(\Equal6~0_combout ),
	.cout());
defparam \Equal6~0 .lut_mask = 16'h00AA;
defparam \Equal6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_num_lines[1]~0 (
	.dataa(\Equal10~0_combout ),
	.datab(\Equal6~0_combout ),
	.datac(gnd),
	.datad(\Equal5~0_combout ),
	.cin(gnd),
	.combout(\addr_num_lines[1]~0_combout ),
	.cout());
defparam \addr_num_lines[1]~0 .lut_mask = 16'hCCAA;
defparam \addr_num_lines[1]~0 .sum_lutc_input = "datac";

dffeas \header_information[18] (
	.clk(clk_clk),
	.d(in_cmd_data[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\header_information[18]~q ),
	.prn(vcc));
defparam \header_information[18] .is_wysiwyg = "true";
defparam \header_information[18] .power_up = "low";

cycloneive_lcell_comb \Add2~0 (
	.dataa(\header_information[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add2~0_combout ),
	.cout(\Add2~1 ));
defparam \Add2~0 .lut_mask = 16'h55AA;
defparam \Add2~0 .sum_lutc_input = "datac";

dffeas \header_information[19] (
	.clk(clk_clk),
	.d(in_cmd_data[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\header_information[19]~q ),
	.prn(vcc));
defparam \header_information[19] .is_wysiwyg = "true";
defparam \header_information[19] .power_up = "low";

cycloneive_lcell_comb \Add2~2 (
	.dataa(\header_information[19]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~1 ),
	.combout(\Add2~2_combout ),
	.cout(\Add2~3 ));
defparam \Add2~2 .lut_mask = 16'hA505;
defparam \Add2~2 .sum_lutc_input = "cin";

cycloneive_lcell_comb \data_in_cnt[0]~8 (
	.dataa(\data_in_cnt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\data_in_cnt[0]~8_combout ),
	.cout(\data_in_cnt[0]~9 ));
defparam \data_in_cnt[0]~8 .lut_mask = 16'h55AA;
defparam \data_in_cnt[0]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb data_in_cnt_done(
	.dataa(Selector8),
	.datab(\data_in_cnt_done~4_combout ),
	.datac(sink_ready),
	.datad(WideOr03),
	.cin(gnd),
	.combout(\data_in_cnt_done~combout ),
	.cout());
defparam data_in_cnt_done.lut_mask = 16'h8880;
defparam data_in_cnt_done.sum_lutc_input = "datac";

cycloneive_lcell_comb \always8~0 (
	.dataa(stateST_SEND_DATA),
	.datab(Selector8),
	.datac(sink_ready),
	.datad(WideOr03),
	.cin(gnd),
	.combout(\always8~0_combout ),
	.cout());
defparam \always8~0 .lut_mask = 16'h8880;
defparam \always8~0 .sum_lutc_input = "datac";

dffeas \data_in_cnt[0] (
	.clk(clk_clk),
	.d(\data_in_cnt[0]~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\data_in_cnt_done~combout ),
	.sload(gnd),
	.ena(\always8~0_combout ),
	.q(\data_in_cnt[0]~q ),
	.prn(vcc));
defparam \data_in_cnt[0] .is_wysiwyg = "true";
defparam \data_in_cnt[0] .power_up = "low";

cycloneive_lcell_comb \data_in_cnt[1]~10 (
	.dataa(\data_in_cnt[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_in_cnt[0]~9 ),
	.combout(\data_in_cnt[1]~10_combout ),
	.cout(\data_in_cnt[1]~11 ));
defparam \data_in_cnt[1]~10 .lut_mask = 16'h5A5F;
defparam \data_in_cnt[1]~10 .sum_lutc_input = "cin";

dffeas \data_in_cnt[1] (
	.clk(clk_clk),
	.d(\data_in_cnt[1]~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\data_in_cnt_done~combout ),
	.sload(gnd),
	.ena(\always8~0_combout ),
	.q(\data_in_cnt[1]~q ),
	.prn(vcc));
defparam \data_in_cnt[1] .is_wysiwyg = "true";
defparam \data_in_cnt[1] .power_up = "low";

cycloneive_lcell_comb \data_in_cnt_done~0 (
	.dataa(\Add2~0_combout ),
	.datab(\Add2~2_combout ),
	.datac(\data_in_cnt[1]~q ),
	.datad(\data_in_cnt[0]~q ),
	.cin(gnd),
	.combout(\data_in_cnt_done~0_combout ),
	.cout());
defparam \data_in_cnt_done~0 .lut_mask = 16'h8241;
defparam \data_in_cnt_done~0 .sum_lutc_input = "datac";

dffeas \header_information[21] (
	.clk(clk_clk),
	.d(in_cmd_data[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\header_information[21]~q ),
	.prn(vcc));
defparam \header_information[21] .is_wysiwyg = "true";
defparam \header_information[21] .power_up = "low";

dffeas \header_information[20] (
	.clk(clk_clk),
	.d(in_cmd_data[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\header_information[20]~q ),
	.prn(vcc));
defparam \header_information[20] .is_wysiwyg = "true";
defparam \header_information[20] .power_up = "low";

cycloneive_lcell_comb \Add2~4 (
	.dataa(\header_information[20]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~3 ),
	.combout(\Add2~4_combout ),
	.cout(\Add2~5 ));
defparam \Add2~4 .lut_mask = 16'h5AAF;
defparam \Add2~4 .sum_lutc_input = "cin";

cycloneive_lcell_comb \Add2~6 (
	.dataa(\header_information[21]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~5 ),
	.combout(\Add2~6_combout ),
	.cout(\Add2~7 ));
defparam \Add2~6 .lut_mask = 16'hA505;
defparam \Add2~6 .sum_lutc_input = "cin";

cycloneive_lcell_comb \data_in_cnt[2]~12 (
	.dataa(\data_in_cnt[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_in_cnt[1]~11 ),
	.combout(\data_in_cnt[2]~12_combout ),
	.cout(\data_in_cnt[2]~13 ));
defparam \data_in_cnt[2]~12 .lut_mask = 16'hA50A;
defparam \data_in_cnt[2]~12 .sum_lutc_input = "cin";

dffeas \data_in_cnt[2] (
	.clk(clk_clk),
	.d(\data_in_cnt[2]~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\data_in_cnt_done~combout ),
	.sload(gnd),
	.ena(\always8~0_combout ),
	.q(\data_in_cnt[2]~q ),
	.prn(vcc));
defparam \data_in_cnt[2] .is_wysiwyg = "true";
defparam \data_in_cnt[2] .power_up = "low";

cycloneive_lcell_comb \data_in_cnt[3]~14 (
	.dataa(\data_in_cnt[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_in_cnt[2]~13 ),
	.combout(\data_in_cnt[3]~14_combout ),
	.cout(\data_in_cnt[3]~15 ));
defparam \data_in_cnt[3]~14 .lut_mask = 16'h5A5F;
defparam \data_in_cnt[3]~14 .sum_lutc_input = "cin";

dffeas \data_in_cnt[3] (
	.clk(clk_clk),
	.d(\data_in_cnt[3]~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\data_in_cnt_done~combout ),
	.sload(gnd),
	.ena(\always8~0_combout ),
	.q(\data_in_cnt[3]~q ),
	.prn(vcc));
defparam \data_in_cnt[3] .is_wysiwyg = "true";
defparam \data_in_cnt[3] .power_up = "low";

cycloneive_lcell_comb \Equal16~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\Add2~4_combout ),
	.datad(\data_in_cnt[2]~q ),
	.cin(gnd),
	.combout(\Equal16~0_combout ),
	.cout());
defparam \Equal16~0 .lut_mask = 16'h0FF0;
defparam \Equal16~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_in_cnt_done~1 (
	.dataa(\data_in_cnt_done~0_combout ),
	.datab(\Add2~6_combout ),
	.datac(\data_in_cnt[3]~q ),
	.datad(\Equal16~0_combout ),
	.cin(gnd),
	.combout(\data_in_cnt_done~1_combout ),
	.cout());
defparam \data_in_cnt_done~1 .lut_mask = 16'h0082;
defparam \data_in_cnt_done~1 .sum_lutc_input = "datac";

dffeas \header_information[22] (
	.clk(clk_clk),
	.d(in_cmd_data[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\header_information[22]~q ),
	.prn(vcc));
defparam \header_information[22] .is_wysiwyg = "true";
defparam \header_information[22] .power_up = "low";

cycloneive_lcell_comb \Add2~8 (
	.dataa(\header_information[22]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~7 ),
	.combout(\Add2~8_combout ),
	.cout(\Add2~9 ));
defparam \Add2~8 .lut_mask = 16'h5AAF;
defparam \Add2~8 .sum_lutc_input = "cin";

dffeas \header_information[23] (
	.clk(clk_clk),
	.d(in_cmd_data[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\header_information[23]~q ),
	.prn(vcc));
defparam \header_information[23] .is_wysiwyg = "true";
defparam \header_information[23] .power_up = "low";

cycloneive_lcell_comb \Add2~10 (
	.dataa(\header_information[23]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~9 ),
	.combout(\Add2~10_combout ),
	.cout(\Add2~11 ));
defparam \Add2~10 .lut_mask = 16'hA505;
defparam \Add2~10 .sum_lutc_input = "cin";

cycloneive_lcell_comb \data_in_cnt[4]~16 (
	.dataa(\data_in_cnt[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_in_cnt[3]~15 ),
	.combout(\data_in_cnt[4]~16_combout ),
	.cout(\data_in_cnt[4]~17 ));
defparam \data_in_cnt[4]~16 .lut_mask = 16'hA50A;
defparam \data_in_cnt[4]~16 .sum_lutc_input = "cin";

dffeas \data_in_cnt[4] (
	.clk(clk_clk),
	.d(\data_in_cnt[4]~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\data_in_cnt_done~combout ),
	.sload(gnd),
	.ena(\always8~0_combout ),
	.q(\data_in_cnt[4]~q ),
	.prn(vcc));
defparam \data_in_cnt[4] .is_wysiwyg = "true";
defparam \data_in_cnt[4] .power_up = "low";

cycloneive_lcell_comb \data_in_cnt[5]~18 (
	.dataa(\data_in_cnt[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_in_cnt[4]~17 ),
	.combout(\data_in_cnt[5]~18_combout ),
	.cout(\data_in_cnt[5]~19 ));
defparam \data_in_cnt[5]~18 .lut_mask = 16'h5A5F;
defparam \data_in_cnt[5]~18 .sum_lutc_input = "cin";

dffeas \data_in_cnt[5] (
	.clk(clk_clk),
	.d(\data_in_cnt[5]~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\data_in_cnt_done~combout ),
	.sload(gnd),
	.ena(\always8~0_combout ),
	.q(\data_in_cnt[5]~q ),
	.prn(vcc));
defparam \data_in_cnt[5] .is_wysiwyg = "true";
defparam \data_in_cnt[5] .power_up = "low";

cycloneive_lcell_comb \data_in_cnt_done~2 (
	.dataa(\Add2~8_combout ),
	.datab(\Add2~10_combout ),
	.datac(\data_in_cnt[5]~q ),
	.datad(\data_in_cnt[4]~q ),
	.cin(gnd),
	.combout(\data_in_cnt_done~2_combout ),
	.cout());
defparam \data_in_cnt_done~2 .lut_mask = 16'h8241;
defparam \data_in_cnt_done~2 .sum_lutc_input = "datac";

dffeas \header_information[24] (
	.clk(clk_clk),
	.d(in_cmd_data[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\header_information[24]~q ),
	.prn(vcc));
defparam \header_information[24] .is_wysiwyg = "true";
defparam \header_information[24] .power_up = "low";

cycloneive_lcell_comb \Add2~12 (
	.dataa(\header_information[24]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~11 ),
	.combout(\Add2~12_combout ),
	.cout(\Add2~13 ));
defparam \Add2~12 .lut_mask = 16'h5AAF;
defparam \Add2~12 .sum_lutc_input = "cin";

dffeas \header_information[25] (
	.clk(clk_clk),
	.d(in_cmd_data[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\header_information[25]~q ),
	.prn(vcc));
defparam \header_information[25] .is_wysiwyg = "true";
defparam \header_information[25] .power_up = "low";

cycloneive_lcell_comb \Add2~14 (
	.dataa(\header_information[25]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~13 ),
	.combout(\Add2~14_combout ),
	.cout(\Add2~15 ));
defparam \Add2~14 .lut_mask = 16'hA505;
defparam \Add2~14 .sum_lutc_input = "cin";

cycloneive_lcell_comb \data_in_cnt[6]~20 (
	.dataa(\data_in_cnt[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_in_cnt[5]~19 ),
	.combout(\data_in_cnt[6]~20_combout ),
	.cout(\data_in_cnt[6]~21 ));
defparam \data_in_cnt[6]~20 .lut_mask = 16'hA50A;
defparam \data_in_cnt[6]~20 .sum_lutc_input = "cin";

dffeas \data_in_cnt[6] (
	.clk(clk_clk),
	.d(\data_in_cnt[6]~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\data_in_cnt_done~combout ),
	.sload(gnd),
	.ena(\always8~0_combout ),
	.q(\data_in_cnt[6]~q ),
	.prn(vcc));
defparam \data_in_cnt[6] .is_wysiwyg = "true";
defparam \data_in_cnt[6] .power_up = "low";

cycloneive_lcell_comb \data_in_cnt[7]~22 (
	.dataa(\data_in_cnt[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\data_in_cnt[6]~21 ),
	.combout(\data_in_cnt[7]~22_combout ),
	.cout());
defparam \data_in_cnt[7]~22 .lut_mask = 16'h5A5A;
defparam \data_in_cnt[7]~22 .sum_lutc_input = "cin";

dffeas \data_in_cnt[7] (
	.clk(clk_clk),
	.d(\data_in_cnt[7]~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\data_in_cnt_done~combout ),
	.sload(gnd),
	.ena(\always8~0_combout ),
	.q(\data_in_cnt[7]~q ),
	.prn(vcc));
defparam \data_in_cnt[7] .is_wysiwyg = "true";
defparam \data_in_cnt[7] .power_up = "low";

cycloneive_lcell_comb \data_in_cnt_done~3 (
	.dataa(\Add2~12_combout ),
	.datab(\Add2~14_combout ),
	.datac(\data_in_cnt[7]~q ),
	.datad(\data_in_cnt[6]~q ),
	.cin(gnd),
	.combout(\data_in_cnt_done~3_combout ),
	.cout());
defparam \data_in_cnt_done~3 .lut_mask = 16'h8241;
defparam \data_in_cnt_done~3 .sum_lutc_input = "datac";

dffeas \header_information[26] (
	.clk(clk_clk),
	.d(in_cmd_data[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\header_information[26]~q ),
	.prn(vcc));
defparam \header_information[26] .is_wysiwyg = "true";
defparam \header_information[26] .power_up = "low";

cycloneive_lcell_comb \Add2~16 (
	.dataa(\header_information[26]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add2~15 ),
	.combout(\Add2~16_combout ),
	.cout());
defparam \Add2~16 .lut_mask = 16'h5A5A;
defparam \Add2~16 .sum_lutc_input = "cin";

cycloneive_lcell_comb \data_in_cnt_done~4 (
	.dataa(\data_in_cnt_done~1_combout ),
	.datab(\data_in_cnt_done~2_combout ),
	.datac(\data_in_cnt_done~3_combout ),
	.datad(\Add2~16_combout ),
	.cin(gnd),
	.combout(\data_in_cnt_done~4_combout ),
	.cout());
defparam \data_in_cnt_done~4 .lut_mask = 16'h0080;
defparam \data_in_cnt_done~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector5~2 (
	.dataa(\state.ST_WAIT_BUFFER~q ),
	.datab(\buffer_cnt[2]~q ),
	.datac(\buffer_cnt[1]~q ),
	.datad(\buffer_cnt[0]~q ),
	.cin(gnd),
	.combout(\Selector5~2_combout ),
	.cout());
defparam \Selector5~2 .lut_mask = 16'h2AAA;
defparam \Selector5~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector5~3 (
	.dataa(stateST_SEND_DATA),
	.datab(header_information_11),
	.datac(Selector8),
	.datad(\Selector5~2_combout ),
	.cin(gnd),
	.combout(\Selector5~3_combout ),
	.cout());
defparam \Selector5~3 .lut_mask = 16'hFF20;
defparam \Selector5~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector5~7 (
	.dataa(in_ready),
	.datab(demux_channel_2),
	.datac(WideOr03),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector5~7_combout ),
	.cout());
defparam \Selector5~7 .lut_mask = 16'hF8F8;
defparam \Selector5~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector5~4 (
	.dataa(\data_in_cnt_done~4_combout ),
	.datab(\Selector5~2_combout ),
	.datac(\Selector5~3_combout ),
	.datad(\Selector5~7_combout ),
	.cin(gnd),
	.combout(\Selector5~4_combout ),
	.cout());
defparam \Selector5~4 .lut_mask = 16'hECCC;
defparam \Selector5~4 .sum_lutc_input = "datac";

dffeas \header_information[10] (
	.clk(clk_clk),
	.d(in_cmd_data[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\header_information[10]~q ),
	.prn(vcc));
defparam \header_information[10] .is_wysiwyg = "true";
defparam \header_information[10] .power_up = "low";

cycloneive_lcell_comb \Selector5~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(header_information_11),
	.datad(\header_information[10]~q ),
	.cin(gnd),
	.combout(\Selector5~5_combout ),
	.cout());
defparam \Selector5~5 .lut_mask = 16'h000F;
defparam \Selector5~5 .sum_lutc_input = "datac";

dffeas \header_information[8] (
	.clk(clk_clk),
	.d(in_cmd_data[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\header_information[8]~q ),
	.prn(vcc));
defparam \header_information[8] .is_wysiwyg = "true";
defparam \header_information[8] .power_up = "low";

cycloneive_lcell_comb \Selector3~2 (
	.dataa(stateST_SEND_OPCODE),
	.datab(sink_ready),
	.datac(WideOr03),
	.datad(\header_information[8]~q ),
	.cin(gnd),
	.combout(\Selector3~2_combout ),
	.cout());
defparam \Selector3~2 .lut_mask = 16'h00A8;
defparam \Selector3~2 .sum_lutc_input = "datac";

dffeas \header_information[9] (
	.clk(clk_clk),
	.d(in_cmd_data[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\header_information[9]~q ),
	.prn(vcc));
defparam \header_information[9] .is_wysiwyg = "true";
defparam \header_information[9] .power_up = "low";

cycloneive_lcell_comb \addr_cnt_done~0 (
	.dataa(Selector8),
	.datab(WideOr03),
	.datac(in_ready),
	.datad(demux_channel_2),
	.cin(gnd),
	.combout(\addr_cnt_done~0_combout ),
	.cout());
defparam \addr_cnt_done~0 .lut_mask = 16'hA888;
defparam \addr_cnt_done~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_cnt_next[0]~1 (
	.dataa(\addr_cnt[1]~q ),
	.datab(\header_information[9]~q ),
	.datac(\addr_cnt_done~0_combout ),
	.datad(\addr_cnt[0]~q ),
	.cin(gnd),
	.combout(\addr_cnt_next[0]~1_combout ),
	.cout());
defparam \addr_cnt_next[0]~1 .lut_mask = 16'h00EF;
defparam \addr_cnt_next[0]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_cnt_next[0]~2 (
	.dataa(\addr_cnt_next[0]~1_combout ),
	.datab(\addr_cnt[0]~q ),
	.datac(stateST_SEND_ADDR),
	.datad(WideOr06),
	.cin(gnd),
	.combout(\addr_cnt_next[0]~2_combout ),
	.cout());
defparam \addr_cnt_next[0]~2 .lut_mask = 16'hACCC;
defparam \addr_cnt_next[0]~2 .sum_lutc_input = "datac";

dffeas \addr_cnt[0] (
	.clk(clk_clk),
	.d(\addr_cnt_next[0]~2_combout ),
	.asdata(\header_information[9]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(stateST_SEND_OPCODE),
	.ena(vcc),
	.q(\addr_cnt[0]~q ),
	.prn(vcc));
defparam \addr_cnt[0] .is_wysiwyg = "true";
defparam \addr_cnt[0] .power_up = "low";

cycloneive_lcell_comb \addr_cnt_next[1]~0 (
	.dataa(\addr_cnt[1]~q ),
	.datab(\addr_cnt[0]~q ),
	.datac(stateST_SEND_ADDR),
	.datad(WideOr06),
	.cin(gnd),
	.combout(\addr_cnt_next[1]~0_combout ),
	.cout());
defparam \addr_cnt_next[1]~0 .lut_mask = 16'h9AAA;
defparam \addr_cnt_next[1]~0 .sum_lutc_input = "datac";

dffeas \addr_cnt[1] (
	.clk(clk_clk),
	.d(\addr_cnt_next[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(stateST_SEND_OPCODE),
	.ena(vcc),
	.q(\addr_cnt[1]~q ),
	.prn(vcc));
defparam \addr_cnt[1] .is_wysiwyg = "true";
defparam \addr_cnt[1] .power_up = "low";

cycloneive_lcell_comb \Selector20~0 (
	.dataa(stateST_SEND_ADDR),
	.datab(\addr_cnt[1]~q ),
	.datac(\addr_cnt[0]~q ),
	.datad(Selector8),
	.cin(gnd),
	.combout(\Selector20~0_combout ),
	.cout());
defparam \Selector20~0 .lut_mask = 16'h0200;
defparam \Selector20~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector20~1 (
	.dataa(WideOr03),
	.datab(in_ready),
	.datac(demux_channel_2),
	.datad(\Selector20~0_combout ),
	.cin(gnd),
	.combout(\Selector20~1_combout ),
	.cout());
defparam \Selector20~1 .lut_mask = 16'hEA00;
defparam \Selector20~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector5~6 (
	.dataa(\Selector5~4_combout ),
	.datab(\Selector5~5_combout ),
	.datac(\Selector3~2_combout ),
	.datad(\Selector20~1_combout ),
	.cin(gnd),
	.combout(\Selector5~6_combout ),
	.cout());
defparam \Selector5~6 .lut_mask = 16'hEEEA;
defparam \Selector5~6 .sum_lutc_input = "datac";

dffeas \state.ST_WAIT_BUFFER (
	.clk(clk_clk),
	.d(\Selector5~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_WAIT_BUFFER~q ),
	.prn(vcc));
defparam \state.ST_WAIT_BUFFER .is_wysiwyg = "true";
defparam \state.ST_WAIT_BUFFER .power_up = "low";

cycloneive_lcell_comb \buffer_cnt[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\buffer_cnt[0]~q ),
	.datad(\state.ST_WAIT_BUFFER~q ),
	.cin(gnd),
	.combout(\buffer_cnt[0]~2_combout ),
	.cout());
defparam \buffer_cnt[0]~2 .lut_mask = 16'h0FF0;
defparam \buffer_cnt[0]~2 .sum_lutc_input = "datac";

dffeas \buffer_cnt[0] (
	.clk(clk_clk),
	.d(\buffer_cnt[0]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\buffer_cnt[0]~q ),
	.prn(vcc));
defparam \buffer_cnt[0] .is_wysiwyg = "true";
defparam \buffer_cnt[0] .power_up = "low";

cycloneive_lcell_comb \buffer_cnt[1]~1 (
	.dataa(gnd),
	.datab(\buffer_cnt[1]~q ),
	.datac(\buffer_cnt[0]~q ),
	.datad(\state.ST_WAIT_BUFFER~q ),
	.cin(gnd),
	.combout(\buffer_cnt[1]~1_combout ),
	.cout());
defparam \buffer_cnt[1]~1 .lut_mask = 16'h3CCC;
defparam \buffer_cnt[1]~1 .sum_lutc_input = "datac";

dffeas \buffer_cnt[1] (
	.clk(clk_clk),
	.d(\buffer_cnt[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\buffer_cnt[1]~q ),
	.prn(vcc));
defparam \buffer_cnt[1] .is_wysiwyg = "true";
defparam \buffer_cnt[1] .power_up = "low";

cycloneive_lcell_comb \buffer_cnt[2]~0 (
	.dataa(\buffer_cnt[2]~q ),
	.datab(\buffer_cnt[1]~q ),
	.datac(\buffer_cnt[0]~q ),
	.datad(\state.ST_WAIT_BUFFER~q ),
	.cin(gnd),
	.combout(\buffer_cnt[2]~0_combout ),
	.cout());
defparam \buffer_cnt[2]~0 .lut_mask = 16'h6AAA;
defparam \buffer_cnt[2]~0 .sum_lutc_input = "datac";

dffeas \buffer_cnt[2] (
	.clk(clk_clk),
	.d(\buffer_cnt[2]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\buffer_cnt[2]~q ),
	.prn(vcc));
defparam \buffer_cnt[2] .is_wysiwyg = "true";
defparam \buffer_cnt[2] .power_up = "low";

cycloneive_lcell_comb \Selector6~0 (
	.dataa(\buffer_cnt[2]~q ),
	.datab(\buffer_cnt[1]~q ),
	.datac(\buffer_cnt[0]~q ),
	.datad(\state.ST_WAIT_BUFFER~q ),
	.cin(gnd),
	.combout(\Selector6~0_combout ),
	.cout());
defparam \Selector6~0 .lut_mask = 16'h8000;
defparam \Selector6~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector6~1 (
	.dataa(\Selector6~0_combout ),
	.datab(stateST_SEND_DUMMY_RSP),
	.datac(gnd),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\Selector6~1_combout ),
	.cout());
defparam \Selector6~1 .lut_mask = 16'hAAEE;
defparam \Selector6~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_out_cnt[0]~8 (
	.dataa(\data_out_cnt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\data_out_cnt[0]~8_combout ),
	.cout(\data_out_cnt[0]~9 ));
defparam \data_out_cnt[0]~8 .lut_mask = 16'h55AA;
defparam \data_out_cnt[0]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \always12~1 (
	.dataa(out_rsp_valid),
	.datab(\state.ST_WAIT_RSP~q ),
	.datac(\data_adapter_8_32_inst|a_ready~combout ),
	.datad(\data_adapter_8_32_inst|a_valid~q ),
	.cin(gnd),
	.combout(\always12~1_combout ),
	.cout());
defparam \always12~1 .lut_mask = 16'h8088;
defparam \always12~1 .sum_lutc_input = "datac";

dffeas \data_out_cnt[0] (
	.clk(clk_clk),
	.d(\data_out_cnt[0]~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\in_rsp_eop~combout ),
	.sload(gnd),
	.ena(\always12~1_combout ),
	.q(\data_out_cnt[0]~q ),
	.prn(vcc));
defparam \data_out_cnt[0] .is_wysiwyg = "true";
defparam \data_out_cnt[0] .power_up = "low";

cycloneive_lcell_comb \data_out_cnt[1]~10 (
	.dataa(\data_out_cnt[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_out_cnt[0]~9 ),
	.combout(\data_out_cnt[1]~10_combout ),
	.cout(\data_out_cnt[1]~11 ));
defparam \data_out_cnt[1]~10 .lut_mask = 16'h5A5F;
defparam \data_out_cnt[1]~10 .sum_lutc_input = "cin";

dffeas \data_out_cnt[1] (
	.clk(clk_clk),
	.d(\data_out_cnt[1]~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\in_rsp_eop~combout ),
	.sload(gnd),
	.ena(\always12~1_combout ),
	.q(\data_out_cnt[1]~q ),
	.prn(vcc));
defparam \data_out_cnt[1] .is_wysiwyg = "true";
defparam \data_out_cnt[1] .power_up = "low";

cycloneive_lcell_comb \data_out_cnt[2]~12 (
	.dataa(\data_out_cnt[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_out_cnt[1]~11 ),
	.combout(\data_out_cnt[2]~12_combout ),
	.cout(\data_out_cnt[2]~13 ));
defparam \data_out_cnt[2]~12 .lut_mask = 16'hA50A;
defparam \data_out_cnt[2]~12 .sum_lutc_input = "cin";

dffeas \data_out_cnt[2] (
	.clk(clk_clk),
	.d(\data_out_cnt[2]~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\in_rsp_eop~combout ),
	.sload(gnd),
	.ena(\always12~1_combout ),
	.q(\data_out_cnt[2]~q ),
	.prn(vcc));
defparam \data_out_cnt[2] .is_wysiwyg = "true";
defparam \data_out_cnt[2] .power_up = "low";

cycloneive_lcell_comb \data_out_cnt[3]~14 (
	.dataa(\data_out_cnt[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_out_cnt[2]~13 ),
	.combout(\data_out_cnt[3]~14_combout ),
	.cout(\data_out_cnt[3]~15 ));
defparam \data_out_cnt[3]~14 .lut_mask = 16'h5A5F;
defparam \data_out_cnt[3]~14 .sum_lutc_input = "cin";

dffeas \data_out_cnt[3] (
	.clk(clk_clk),
	.d(\data_out_cnt[3]~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\in_rsp_eop~combout ),
	.sload(gnd),
	.ena(\always12~1_combout ),
	.q(\data_out_cnt[3]~q ),
	.prn(vcc));
defparam \data_out_cnt[3] .is_wysiwyg = "true";
defparam \data_out_cnt[3] .power_up = "low";

cycloneive_lcell_comb \in_rsp_eop~0 (
	.dataa(\Add2~4_combout ),
	.datab(\Add2~6_combout ),
	.datac(\data_out_cnt[3]~q ),
	.datad(\data_out_cnt[2]~q ),
	.cin(gnd),
	.combout(\in_rsp_eop~0_combout ),
	.cout());
defparam \in_rsp_eop~0 .lut_mask = 16'h8241;
defparam \in_rsp_eop~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_out_cnt[4]~16 (
	.dataa(\data_out_cnt[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_out_cnt[3]~15 ),
	.combout(\data_out_cnt[4]~16_combout ),
	.cout(\data_out_cnt[4]~17 ));
defparam \data_out_cnt[4]~16 .lut_mask = 16'hA50A;
defparam \data_out_cnt[4]~16 .sum_lutc_input = "cin";

dffeas \data_out_cnt[4] (
	.clk(clk_clk),
	.d(\data_out_cnt[4]~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\in_rsp_eop~combout ),
	.sload(gnd),
	.ena(\always12~1_combout ),
	.q(\data_out_cnt[4]~q ),
	.prn(vcc));
defparam \data_out_cnt[4] .is_wysiwyg = "true";
defparam \data_out_cnt[4] .power_up = "low";

cycloneive_lcell_comb \data_out_cnt[5]~18 (
	.dataa(\data_out_cnt[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_out_cnt[4]~17 ),
	.combout(\data_out_cnt[5]~18_combout ),
	.cout(\data_out_cnt[5]~19 ));
defparam \data_out_cnt[5]~18 .lut_mask = 16'h5A5F;
defparam \data_out_cnt[5]~18 .sum_lutc_input = "cin";

dffeas \data_out_cnt[5] (
	.clk(clk_clk),
	.d(\data_out_cnt[5]~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\in_rsp_eop~combout ),
	.sload(gnd),
	.ena(\always12~1_combout ),
	.q(\data_out_cnt[5]~q ),
	.prn(vcc));
defparam \data_out_cnt[5] .is_wysiwyg = "true";
defparam \data_out_cnt[5] .power_up = "low";

cycloneive_lcell_comb \data_out_cnt[6]~20 (
	.dataa(\data_out_cnt[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\data_out_cnt[5]~19 ),
	.combout(\data_out_cnt[6]~20_combout ),
	.cout(\data_out_cnt[6]~21 ));
defparam \data_out_cnt[6]~20 .lut_mask = 16'hA50A;
defparam \data_out_cnt[6]~20 .sum_lutc_input = "cin";

dffeas \data_out_cnt[6] (
	.clk(clk_clk),
	.d(\data_out_cnt[6]~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\in_rsp_eop~combout ),
	.sload(gnd),
	.ena(\always12~1_combout ),
	.q(\data_out_cnt[6]~q ),
	.prn(vcc));
defparam \data_out_cnt[6] .is_wysiwyg = "true";
defparam \data_out_cnt[6] .power_up = "low";

cycloneive_lcell_comb \in_rsp_eop~1 (
	.dataa(\Add2~12_combout ),
	.datab(\data_out_cnt[6]~q ),
	.datac(\Add2~10_combout ),
	.datad(\data_out_cnt[5]~q ),
	.cin(gnd),
	.combout(\in_rsp_eop~1_combout ),
	.cout());
defparam \in_rsp_eop~1 .lut_mask = 16'h9009;
defparam \in_rsp_eop~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \in_rsp_eop~2 (
	.dataa(\Add2~0_combout ),
	.datab(\Add2~2_combout ),
	.datac(\data_out_cnt[1]~q ),
	.datad(\data_out_cnt[0]~q ),
	.cin(gnd),
	.combout(\in_rsp_eop~2_combout ),
	.cout());
defparam \in_rsp_eop~2 .lut_mask = 16'h8241;
defparam \in_rsp_eop~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_out_cnt[7]~22 (
	.dataa(\data_out_cnt[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\data_out_cnt[6]~21 ),
	.combout(\data_out_cnt[7]~22_combout ),
	.cout());
defparam \data_out_cnt[7]~22 .lut_mask = 16'h5A5A;
defparam \data_out_cnt[7]~22 .sum_lutc_input = "cin";

dffeas \data_out_cnt[7] (
	.clk(clk_clk),
	.d(\data_out_cnt[7]~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\in_rsp_eop~combout ),
	.sload(gnd),
	.ena(\always12~1_combout ),
	.q(\data_out_cnt[7]~q ),
	.prn(vcc));
defparam \data_out_cnt[7] .is_wysiwyg = "true";
defparam \data_out_cnt[7] .power_up = "low";

cycloneive_lcell_comb \in_rsp_eop~3 (
	.dataa(\data_adapter_8_32_inst|in_ready~combout ),
	.datab(out_rsp_valid),
	.datac(\Add2~8_combout ),
	.datad(\data_out_cnt[4]~q ),
	.cin(gnd),
	.combout(\in_rsp_eop~3_combout ),
	.cout());
defparam \in_rsp_eop~3 .lut_mask = 16'h8008;
defparam \in_rsp_eop~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \in_rsp_eop~4 (
	.dataa(\in_rsp_eop~2_combout ),
	.datab(\Add2~14_combout ),
	.datac(\data_out_cnt[7]~q ),
	.datad(\in_rsp_eop~3_combout ),
	.cin(gnd),
	.combout(\in_rsp_eop~4_combout ),
	.cout());
defparam \in_rsp_eop~4 .lut_mask = 16'h8200;
defparam \in_rsp_eop~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb in_rsp_eop(
	.dataa(\in_rsp_eop~0_combout ),
	.datab(\Add2~16_combout ),
	.datac(\in_rsp_eop~1_combout ),
	.datad(\in_rsp_eop~4_combout ),
	.cin(gnd),
	.combout(\in_rsp_eop~combout ),
	.cout());
defparam in_rsp_eop.lut_mask = 16'h2000;
defparam in_rsp_eop.sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector4~0 (
	.dataa(stateST_SEND_DATA),
	.datab(\addr_cnt_done~0_combout ),
	.datac(\data_in_cnt_done~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector4~0_combout ),
	.cout());
defparam \Selector4~0 .lut_mask = 16'h8080;
defparam \Selector4~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector4~1 (
	.dataa(\Selector3~2_combout ),
	.datab(\header_information[10]~q ),
	.datac(\Selector20~1_combout ),
	.datad(\Selector4~0_combout ),
	.cin(gnd),
	.combout(\Selector4~1_combout ),
	.cout());
defparam \Selector4~1 .lut_mask = 16'hFF32;
defparam \Selector4~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector4~2 (
	.dataa(\state.ST_WAIT_RSP~q ),
	.datab(\in_rsp_eop~combout ),
	.datac(header_information_11),
	.datad(\Selector4~1_combout ),
	.cin(gnd),
	.combout(\Selector4~2_combout ),
	.cout());
defparam \Selector4~2 .lut_mask = 16'hF222;
defparam \Selector4~2 .sum_lutc_input = "datac";

dffeas \state.ST_WAIT_RSP (
	.clk(clk_clk),
	.d(\Selector4~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_WAIT_RSP~q ),
	.prn(vcc));
defparam \state.ST_WAIT_RSP .is_wysiwyg = "true";
defparam \state.ST_WAIT_RSP .power_up = "low";

cycloneive_lcell_comb \Selector7~0 (
	.dataa(out_valid),
	.datab(out_endofpacket),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector7~0_combout ),
	.cout());
defparam \Selector7~0 .lut_mask = 16'h8888;
defparam \Selector7~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector7~1 (
	.dataa(\state.ST_WAIT_RSP~q ),
	.datab(\in_rsp_eop~combout ),
	.datac(\state.ST_COMPLETE~q ),
	.datad(\Selector7~0_combout ),
	.cin(gnd),
	.combout(\Selector7~1_combout ),
	.cout());
defparam \Selector7~1 .lut_mask = 16'h88F8;
defparam \Selector7~1 .sum_lutc_input = "datac";

dffeas \state.ST_COMPLETE (
	.clk(clk_clk),
	.d(\Selector7~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.ST_COMPLETE~q ),
	.prn(vcc));
defparam \state.ST_COMPLETE .is_wysiwyg = "true";
defparam \state.ST_COMPLETE .power_up = "low";

cycloneive_lcell_comb \Selector0~0 (
	.dataa(stateST_SEND_DUMMY_RSP),
	.datab(\state.ST_COMPLETE~q ),
	.datac(\Selector7~0_combout ),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
defparam \Selector0~0 .lut_mask = 16'hEAC8;
defparam \Selector0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector0~1 (
	.dataa(\Selector0~0_combout ),
	.datab(WideOr1),
	.datac(src_startofpacket),
	.datad(stateST_IDLE),
	.cin(gnd),
	.combout(\Selector0~1_combout ),
	.cout());
defparam \Selector0~1 .lut_mask = 16'h5540;
defparam \Selector0~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector3~6 (
	.dataa(in_ready),
	.datab(demux_channel_2),
	.datac(WideOr03),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector3~6_combout ),
	.cout());
defparam \Selector3~6 .lut_mask = 16'h0707;
defparam \Selector3~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector3~3 (
	.dataa(stateST_SEND_DATA),
	.datab(Selector8),
	.datac(\data_in_cnt_done~4_combout ),
	.datad(\Selector3~6_combout ),
	.cin(gnd),
	.combout(\Selector3~3_combout ),
	.cout());
defparam \Selector3~3 .lut_mask = 16'hAA2A;
defparam \Selector3~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector3~4 (
	.dataa(\Selector3~3_combout ),
	.datab(\header_information[10]~q ),
	.datac(\Selector3~2_combout ),
	.datad(\Selector20~1_combout ),
	.cin(gnd),
	.combout(\Selector3~4_combout ),
	.cout());
defparam \Selector3~4 .lut_mask = 16'hEEEA;
defparam \Selector3~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~0 (
	.dataa(WideOr05),
	.datab(in_ready),
	.datac(op_num_lines_2),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
defparam \Selector2~0 .lut_mask = 16'hEAEA;
defparam \Selector2~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~1 (
	.dataa(\addr_cnt[1]~q ),
	.datab(\addr_cnt[0]~q ),
	.datac(stateST_SEND_ADDR),
	.datad(WideOr06),
	.cin(gnd),
	.combout(\Selector2~1_combout ),
	.cout());
defparam \Selector2~1 .lut_mask = 16'hE0F0;
defparam \Selector2~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector2~2 (
	.dataa(\header_information[8]~q ),
	.datab(stateST_SEND_OPCODE),
	.datac(\Selector2~0_combout ),
	.datad(\Selector2~1_combout ),
	.cin(gnd),
	.combout(\Selector2~2_combout ),
	.cout());
defparam \Selector2~2 .lut_mask = 16'hFF80;
defparam \Selector2~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector18~0 (
	.dataa(\data_adapter_32_8_inst|state_register[1]~q ),
	.datab(\data_adapter_32_8_inst|state_register[0]~q ),
	.datac(\data_adapter_32_8_inst|out_valid~q ),
	.datad(\data_adapter_32_8_inst|a_valid~q ),
	.cin(gnd),
	.combout(\Selector18~0_combout ),
	.cout());
defparam \Selector18~0 .lut_mask = 16'h08FF;
defparam \Selector18~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \last_word_detect~0 (
	.dataa(\Selector5~5_combout ),
	.datab(src_payload_0),
	.datac(WideOr1),
	.datad(Selector182),
	.cin(gnd),
	.combout(\last_word_detect~0_combout ),
	.cout());
defparam \last_word_detect~0 .lut_mask = 16'h4000;
defparam \last_word_detect~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \last_word_detect~1 (
	.dataa(\last_word_detect~q ),
	.datab(stateST_SEND_DUMMY_RSP),
	.datac(\state.ST_COMPLETE~q ),
	.datad(\last_word_detect~0_combout ),
	.cin(gnd),
	.combout(\last_word_detect~1_combout ),
	.cout());
defparam \last_word_detect~1 .lut_mask = 16'h0302;
defparam \last_word_detect~1 .sum_lutc_input = "datac";

dffeas last_word_detect(
	.clk(clk_clk),
	.d(\last_word_detect~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset),
	.sload(gnd),
	.ena(vcc),
	.q(\last_word_detect~q ),
	.prn(vcc));
defparam last_word_detect.is_wysiwyg = "true";
defparam last_word_detect.power_up = "low";

cycloneive_lcell_comb \Selector18~1 (
	.dataa(stateST_SEND_DATA),
	.datab(stateST_SEND_ADDR),
	.datac(gnd),
	.datad(\last_word_detect~q ),
	.cin(gnd),
	.combout(\Selector18~1_combout ),
	.cout());
defparam \Selector18~1 .lut_mask = 16'h00EE;
defparam \Selector18~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_num_lines~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(csr_op_protocol_data_8),
	.datad(csr_op_protocol_data_9),
	.cin(gnd),
	.combout(\data_num_lines~5_combout ),
	.cout());
defparam \data_num_lines~5 .lut_mask = 16'h0FF0;
defparam \data_num_lines~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_num_lines~6 (
	.dataa(\data_num_lines~5_combout ),
	.datab(\Equal5~0_combout ),
	.datac(csr_op_protocol_data_16),
	.datad(csr_op_protocol_data_17),
	.cin(gnd),
	.combout(\data_num_lines~6_combout ),
	.cout());
defparam \data_num_lines~6 .lut_mask = 16'h8BB8;
defparam \data_num_lines~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_num_lines~9 (
	.dataa(csr_op_protocol_data_0),
	.datab(csr_op_protocol_data_1),
	.datac(\data_num_lines~6_combout ),
	.datad(\always2~1_combout ),
	.cin(gnd),
	.combout(\data_num_lines~9_combout ),
	.cout());
defparam \data_num_lines~9 .lut_mask = 16'h990F;
defparam \data_num_lines~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data_num_lines~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(csr_op_protocol_data_0),
	.datad(csr_op_protocol_data_1),
	.cin(gnd),
	.combout(\data_num_lines~4_combout ),
	.cout());
defparam \data_num_lines~4 .lut_mask = 16'hF00F;
defparam \data_num_lines~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector18~4 (
	.dataa(in_ready),
	.datab(WideOr02),
	.datac(WideOr01),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector18~4_combout ),
	.cout());
defparam \Selector18~4 .lut_mask = 16'hF8F8;
defparam \Selector18~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector1~0 (
	.dataa(\always0~0_combout ),
	.datab(stateST_SEND_OPCODE),
	.datac(stateST_IDLE),
	.datad(WideOr07),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'h0ACE;
defparam \Selector1~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_num_lines~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(csr_op_protocol_data_4),
	.datad(csr_op_protocol_data_5),
	.cin(gnd),
	.combout(\addr_num_lines~6_combout ),
	.cout());
defparam \addr_num_lines~6 .lut_mask = 16'h0FF0;
defparam \addr_num_lines~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_num_lines~7 (
	.dataa(\addr_num_lines~6_combout ),
	.datab(\Equal5~0_combout ),
	.datac(csr_op_protocol_data_12),
	.datad(csr_op_protocol_data_13),
	.cin(gnd),
	.combout(\addr_num_lines~7_combout ),
	.cout());
defparam \addr_num_lines~7 .lut_mask = 16'h8BB8;
defparam \addr_num_lines~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_num_lines~8 (
	.dataa(csr_op_protocol_data_0),
	.datab(csr_op_protocol_data_1),
	.datac(\addr_num_lines~7_combout ),
	.datad(\always2~1_combout ),
	.cin(gnd),
	.combout(\addr_num_lines~8_combout ),
	.cout());
defparam \addr_num_lines~8 .lut_mask = 16'h990F;
defparam \addr_num_lines~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal0~0 (
	.dataa(in_cmd_channel[1]),
	.datab(gnd),
	.datac(gnd),
	.datad(in_cmd_channel[0]),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h00AA;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_mem~0 (
	.dataa(csr_flash_cmd_addr_data_8),
	.datab(has_addr),
	.datac(mem_addr_reg_6),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\addr_mem~0_combout ),
	.cout());
defparam \addr_mem~0 .lut_mask = 16'h88F0;
defparam \addr_mem~0 .sum_lutc_input = "datac";

dffeas \addr_mem[1][0] (
	.clk(clk_clk),
	.d(\addr_mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[1][0]~q ),
	.prn(vcc));
defparam \addr_mem[1][0] .is_wysiwyg = "true";
defparam \addr_mem[1][0] .power_up = "low";

cycloneive_lcell_comb \addr_mem~1 (
	.dataa(csr_flash_cmd_addr_data_16),
	.datab(has_addr),
	.datac(mem_addr_reg_14),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\addr_mem~1_combout ),
	.cout());
defparam \addr_mem~1 .lut_mask = 16'h88F0;
defparam \addr_mem~1 .sum_lutc_input = "datac";

dffeas \addr_mem[2][0] (
	.clk(clk_clk),
	.d(\addr_mem~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[2][0]~q ),
	.prn(vcc));
defparam \addr_mem[2][0] .is_wysiwyg = "true";
defparam \addr_mem[2][0] .power_up = "low";

cycloneive_lcell_comb \addr_mem~2 (
	.dataa(csr_flash_cmd_addr_data_0),
	.datab(has_addr),
	.datac(addr_bytes_xip_0),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\addr_mem~2_combout ),
	.cout());
defparam \addr_mem~2 .lut_mask = 16'h88F0;
defparam \addr_mem~2 .sum_lutc_input = "datac";

dffeas \addr_mem[0][0] (
	.clk(clk_clk),
	.d(\addr_mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[0][0]~q ),
	.prn(vcc));
defparam \addr_mem[0][0] .is_wysiwyg = "true";
defparam \addr_mem[0][0] .power_up = "low";

cycloneive_lcell_comb \Selector16~0 (
	.dataa(\addr_cnt[0]~q ),
	.datab(\addr_mem[2][0]~q ),
	.datac(\addr_cnt[1]~q ),
	.datad(\addr_mem[0][0]~q ),
	.cin(gnd),
	.combout(\Selector16~0_combout ),
	.cout());
defparam \Selector16~0 .lut_mask = 16'hE5E0;
defparam \Selector16~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_mem~3 (
	.dataa(csr_flash_cmd_addr_data_24),
	.datab(in_cmd_channel[1]),
	.datac(has_addr),
	.datad(in_cmd_channel[0]),
	.cin(gnd),
	.combout(\addr_mem~3_combout ),
	.cout());
defparam \addr_mem~3 .lut_mask = 16'h0080;
defparam \addr_mem~3 .sum_lutc_input = "datac";

dffeas \addr_mem[3][0] (
	.clk(clk_clk),
	.d(\addr_mem~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[3][0]~q ),
	.prn(vcc));
defparam \addr_mem[3][0] .is_wysiwyg = "true";
defparam \addr_mem[3][0] .power_up = "low";

cycloneive_lcell_comb \Selector16~1 (
	.dataa(\addr_mem[1][0]~q ),
	.datab(\addr_cnt[0]~q ),
	.datac(\Selector16~0_combout ),
	.datad(\addr_mem[3][0]~q ),
	.cin(gnd),
	.combout(\Selector16~1_combout ),
	.cout());
defparam \Selector16~1 .lut_mask = 16'hF838;
defparam \Selector16~1 .sum_lutc_input = "datac";

dffeas \header_information[0] (
	.clk(clk_clk),
	.d(in_cmd_data[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\header_information[0]~q ),
	.prn(vcc));
defparam \header_information[0] .is_wysiwyg = "true";
defparam \header_information[0] .power_up = "low";

cycloneive_lcell_comb \Selector16~2 (
	.dataa(\Selector16~1_combout ),
	.datab(stateST_SEND_OPCODE),
	.datac(\header_information[0]~q ),
	.datad(stateST_SEND_ADDR),
	.cin(gnd),
	.combout(\Selector16~2_combout ),
	.cout());
defparam \Selector16~2 .lut_mask = 16'hAAC0;
defparam \Selector16~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_mem~4 (
	.dataa(csr_flash_cmd_addr_data_12),
	.datab(has_addr),
	.datac(mem_addr_reg_10),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\addr_mem~4_combout ),
	.cout());
defparam \addr_mem~4 .lut_mask = 16'h88F0;
defparam \addr_mem~4 .sum_lutc_input = "datac";

dffeas \addr_mem[1][4] (
	.clk(clk_clk),
	.d(\addr_mem~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[1][4]~q ),
	.prn(vcc));
defparam \addr_mem[1][4] .is_wysiwyg = "true";
defparam \addr_mem[1][4] .power_up = "low";

cycloneive_lcell_comb \addr_mem~5 (
	.dataa(csr_flash_cmd_addr_data_20),
	.datab(has_addr),
	.datac(mem_addr_reg_18),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\addr_mem~5_combout ),
	.cout());
defparam \addr_mem~5 .lut_mask = 16'h88F0;
defparam \addr_mem~5 .sum_lutc_input = "datac";

dffeas \addr_mem[2][4] (
	.clk(clk_clk),
	.d(\addr_mem~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[2][4]~q ),
	.prn(vcc));
defparam \addr_mem[2][4] .is_wysiwyg = "true";
defparam \addr_mem[2][4] .power_up = "low";

cycloneive_lcell_comb \addr_mem~6 (
	.dataa(csr_flash_cmd_addr_data_4),
	.datab(has_addr),
	.datac(mem_addr_reg_2),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\addr_mem~6_combout ),
	.cout());
defparam \addr_mem~6 .lut_mask = 16'h88F0;
defparam \addr_mem~6 .sum_lutc_input = "datac";

dffeas \addr_mem[0][4] (
	.clk(clk_clk),
	.d(\addr_mem~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[0][4]~q ),
	.prn(vcc));
defparam \addr_mem[0][4] .is_wysiwyg = "true";
defparam \addr_mem[0][4] .power_up = "low";

cycloneive_lcell_comb \Selector12~0 (
	.dataa(\addr_cnt[0]~q ),
	.datab(\addr_mem[2][4]~q ),
	.datac(\addr_cnt[1]~q ),
	.datad(\addr_mem[0][4]~q ),
	.cin(gnd),
	.combout(\Selector12~0_combout ),
	.cout());
defparam \Selector12~0 .lut_mask = 16'hE5E0;
defparam \Selector12~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_mem~7 (
	.dataa(csr_flash_cmd_addr_data_28),
	.datab(in_cmd_channel[1]),
	.datac(has_addr),
	.datad(in_cmd_channel[0]),
	.cin(gnd),
	.combout(\addr_mem~7_combout ),
	.cout());
defparam \addr_mem~7 .lut_mask = 16'h0080;
defparam \addr_mem~7 .sum_lutc_input = "datac";

dffeas \addr_mem[3][4] (
	.clk(clk_clk),
	.d(\addr_mem~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[3][4]~q ),
	.prn(vcc));
defparam \addr_mem[3][4] .is_wysiwyg = "true";
defparam \addr_mem[3][4] .power_up = "low";

cycloneive_lcell_comb \Selector12~1 (
	.dataa(\addr_mem[1][4]~q ),
	.datab(\addr_cnt[0]~q ),
	.datac(\Selector12~0_combout ),
	.datad(\addr_mem[3][4]~q ),
	.cin(gnd),
	.combout(\Selector12~1_combout ),
	.cout());
defparam \Selector12~1 .lut_mask = 16'hF838;
defparam \Selector12~1 .sum_lutc_input = "datac";

dffeas \header_information[4] (
	.clk(clk_clk),
	.d(in_cmd_data[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\header_information[4]~q ),
	.prn(vcc));
defparam \header_information[4] .is_wysiwyg = "true";
defparam \header_information[4] .power_up = "low";

cycloneive_lcell_comb \Selector12~2 (
	.dataa(\Selector12~1_combout ),
	.datab(stateST_SEND_OPCODE),
	.datac(\header_information[4]~q ),
	.datad(stateST_SEND_ADDR),
	.cin(gnd),
	.combout(\Selector12~2_combout ),
	.cout());
defparam \Selector12~2 .lut_mask = 16'hAAC0;
defparam \Selector12~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_mem~8 (
	.dataa(csr_flash_cmd_addr_data_10),
	.datab(has_addr),
	.datac(mem_addr_reg_8),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\addr_mem~8_combout ),
	.cout());
defparam \addr_mem~8 .lut_mask = 16'h88F0;
defparam \addr_mem~8 .sum_lutc_input = "datac";

dffeas \addr_mem[1][2] (
	.clk(clk_clk),
	.d(\addr_mem~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[1][2]~q ),
	.prn(vcc));
defparam \addr_mem[1][2] .is_wysiwyg = "true";
defparam \addr_mem[1][2] .power_up = "low";

cycloneive_lcell_comb \addr_mem~9 (
	.dataa(csr_flash_cmd_addr_data_18),
	.datab(has_addr),
	.datac(mem_addr_reg_16),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\addr_mem~9_combout ),
	.cout());
defparam \addr_mem~9 .lut_mask = 16'h88F0;
defparam \addr_mem~9 .sum_lutc_input = "datac";

dffeas \addr_mem[2][2] (
	.clk(clk_clk),
	.d(\addr_mem~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[2][2]~q ),
	.prn(vcc));
defparam \addr_mem[2][2] .is_wysiwyg = "true";
defparam \addr_mem[2][2] .power_up = "low";

cycloneive_lcell_comb \addr_mem~10 (
	.dataa(csr_flash_cmd_addr_data_2),
	.datab(has_addr),
	.datac(mem_addr_reg_0),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\addr_mem~10_combout ),
	.cout());
defparam \addr_mem~10 .lut_mask = 16'h88F0;
defparam \addr_mem~10 .sum_lutc_input = "datac";

dffeas \addr_mem[0][2] (
	.clk(clk_clk),
	.d(\addr_mem~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[0][2]~q ),
	.prn(vcc));
defparam \addr_mem[0][2] .is_wysiwyg = "true";
defparam \addr_mem[0][2] .power_up = "low";

cycloneive_lcell_comb \Selector14~0 (
	.dataa(\addr_cnt[0]~q ),
	.datab(\addr_mem[2][2]~q ),
	.datac(\addr_cnt[1]~q ),
	.datad(\addr_mem[0][2]~q ),
	.cin(gnd),
	.combout(\Selector14~0_combout ),
	.cout());
defparam \Selector14~0 .lut_mask = 16'hE5E0;
defparam \Selector14~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_mem~11 (
	.dataa(csr_flash_cmd_addr_data_26),
	.datab(in_cmd_channel[1]),
	.datac(has_addr),
	.datad(in_cmd_channel[0]),
	.cin(gnd),
	.combout(\addr_mem~11_combout ),
	.cout());
defparam \addr_mem~11 .lut_mask = 16'h0080;
defparam \addr_mem~11 .sum_lutc_input = "datac";

dffeas \addr_mem[3][2] (
	.clk(clk_clk),
	.d(\addr_mem~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[3][2]~q ),
	.prn(vcc));
defparam \addr_mem[3][2] .is_wysiwyg = "true";
defparam \addr_mem[3][2] .power_up = "low";

cycloneive_lcell_comb \Selector14~1 (
	.dataa(\addr_mem[1][2]~q ),
	.datab(\addr_cnt[0]~q ),
	.datac(\Selector14~0_combout ),
	.datad(\addr_mem[3][2]~q ),
	.cin(gnd),
	.combout(\Selector14~1_combout ),
	.cout());
defparam \Selector14~1 .lut_mask = 16'hF838;
defparam \Selector14~1 .sum_lutc_input = "datac";

dffeas \header_information[2] (
	.clk(clk_clk),
	.d(in_cmd_data[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\header_information[2]~q ),
	.prn(vcc));
defparam \header_information[2] .is_wysiwyg = "true";
defparam \header_information[2] .power_up = "low";

cycloneive_lcell_comb \Selector14~2 (
	.dataa(\Selector14~1_combout ),
	.datab(stateST_SEND_OPCODE),
	.datac(\header_information[2]~q ),
	.datad(stateST_SEND_ADDR),
	.cin(gnd),
	.combout(\Selector14~2_combout ),
	.cout());
defparam \Selector14~2 .lut_mask = 16'hAAC0;
defparam \Selector14~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_mem~12 (
	.dataa(csr_flash_cmd_addr_data_17),
	.datab(has_addr),
	.datac(mem_addr_reg_15),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\addr_mem~12_combout ),
	.cout());
defparam \addr_mem~12 .lut_mask = 16'h88F0;
defparam \addr_mem~12 .sum_lutc_input = "datac";

dffeas \addr_mem[2][1] (
	.clk(clk_clk),
	.d(\addr_mem~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[2][1]~q ),
	.prn(vcc));
defparam \addr_mem[2][1] .is_wysiwyg = "true";
defparam \addr_mem[2][1] .power_up = "low";

cycloneive_lcell_comb \addr_mem~13 (
	.dataa(csr_flash_cmd_addr_data_9),
	.datab(has_addr),
	.datac(mem_addr_reg_7),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\addr_mem~13_combout ),
	.cout());
defparam \addr_mem~13 .lut_mask = 16'h88F0;
defparam \addr_mem~13 .sum_lutc_input = "datac";

dffeas \addr_mem[1][1] (
	.clk(clk_clk),
	.d(\addr_mem~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[1][1]~q ),
	.prn(vcc));
defparam \addr_mem[1][1] .is_wysiwyg = "true";
defparam \addr_mem[1][1] .power_up = "low";

cycloneive_lcell_comb \addr_mem~14 (
	.dataa(csr_flash_cmd_addr_data_1),
	.datab(has_addr),
	.datac(WideOr19),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\addr_mem~14_combout ),
	.cout());
defparam \addr_mem~14 .lut_mask = 16'h88F0;
defparam \addr_mem~14 .sum_lutc_input = "datac";

dffeas \addr_mem[0][1] (
	.clk(clk_clk),
	.d(\addr_mem~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[0][1]~q ),
	.prn(vcc));
defparam \addr_mem[0][1] .is_wysiwyg = "true";
defparam \addr_mem[0][1] .power_up = "low";

cycloneive_lcell_comb \Selector15~0 (
	.dataa(\addr_cnt[1]~q ),
	.datab(\addr_mem[1][1]~q ),
	.datac(\addr_cnt[0]~q ),
	.datad(\addr_mem[0][1]~q ),
	.cin(gnd),
	.combout(\Selector15~0_combout ),
	.cout());
defparam \Selector15~0 .lut_mask = 16'hE5E0;
defparam \Selector15~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_mem~15 (
	.dataa(csr_flash_cmd_addr_data_25),
	.datab(in_cmd_channel[1]),
	.datac(has_addr),
	.datad(in_cmd_channel[0]),
	.cin(gnd),
	.combout(\addr_mem~15_combout ),
	.cout());
defparam \addr_mem~15 .lut_mask = 16'h0080;
defparam \addr_mem~15 .sum_lutc_input = "datac";

dffeas \addr_mem[3][1] (
	.clk(clk_clk),
	.d(\addr_mem~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[3][1]~q ),
	.prn(vcc));
defparam \addr_mem[3][1] .is_wysiwyg = "true";
defparam \addr_mem[3][1] .power_up = "low";

cycloneive_lcell_comb \Selector15~1 (
	.dataa(\addr_mem[2][1]~q ),
	.datab(\addr_cnt[1]~q ),
	.datac(\Selector15~0_combout ),
	.datad(\addr_mem[3][1]~q ),
	.cin(gnd),
	.combout(\Selector15~1_combout ),
	.cout());
defparam \Selector15~1 .lut_mask = 16'hF838;
defparam \Selector15~1 .sum_lutc_input = "datac";

dffeas \header_information[1] (
	.clk(clk_clk),
	.d(in_cmd_data[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\header_information[1]~q ),
	.prn(vcc));
defparam \header_information[1] .is_wysiwyg = "true";
defparam \header_information[1] .power_up = "low";

cycloneive_lcell_comb \Selector9~0 (
	.dataa(stateST_SEND_DATA),
	.datab(gnd),
	.datac(stateST_SEND_ADDR),
	.datad(stateST_SEND_OPCODE),
	.cin(gnd),
	.combout(\Selector9~0_combout ),
	.cout());
defparam \Selector9~0 .lut_mask = 16'hAAAF;
defparam \Selector9~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector15~2 (
	.dataa(\Selector15~1_combout ),
	.datab(\header_information[1]~q ),
	.datac(stateST_SEND_ADDR),
	.datad(\Selector9~0_combout ),
	.cin(gnd),
	.combout(\Selector15~2_combout ),
	.cout());
defparam \Selector15~2 .lut_mask = 16'h00AC;
defparam \Selector15~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_mem~16 (
	.dataa(csr_flash_cmd_addr_data_19),
	.datab(has_addr),
	.datac(mem_addr_reg_17),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\addr_mem~16_combout ),
	.cout());
defparam \addr_mem~16 .lut_mask = 16'h88F0;
defparam \addr_mem~16 .sum_lutc_input = "datac";

dffeas \addr_mem[2][3] (
	.clk(clk_clk),
	.d(\addr_mem~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[2][3]~q ),
	.prn(vcc));
defparam \addr_mem[2][3] .is_wysiwyg = "true";
defparam \addr_mem[2][3] .power_up = "low";

cycloneive_lcell_comb \addr_mem~17 (
	.dataa(csr_flash_cmd_addr_data_11),
	.datab(has_addr),
	.datac(mem_addr_reg_9),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\addr_mem~17_combout ),
	.cout());
defparam \addr_mem~17 .lut_mask = 16'h88F0;
defparam \addr_mem~17 .sum_lutc_input = "datac";

dffeas \addr_mem[1][3] (
	.clk(clk_clk),
	.d(\addr_mem~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[1][3]~q ),
	.prn(vcc));
defparam \addr_mem[1][3] .is_wysiwyg = "true";
defparam \addr_mem[1][3] .power_up = "low";

cycloneive_lcell_comb \addr_mem~18 (
	.dataa(csr_flash_cmd_addr_data_3),
	.datab(has_addr),
	.datac(mem_addr_reg_1),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\addr_mem~18_combout ),
	.cout());
defparam \addr_mem~18 .lut_mask = 16'h88F0;
defparam \addr_mem~18 .sum_lutc_input = "datac";

dffeas \addr_mem[0][3] (
	.clk(clk_clk),
	.d(\addr_mem~18_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[0][3]~q ),
	.prn(vcc));
defparam \addr_mem[0][3] .is_wysiwyg = "true";
defparam \addr_mem[0][3] .power_up = "low";

cycloneive_lcell_comb \Selector13~0 (
	.dataa(\addr_cnt[1]~q ),
	.datab(\addr_mem[1][3]~q ),
	.datac(\addr_cnt[0]~q ),
	.datad(\addr_mem[0][3]~q ),
	.cin(gnd),
	.combout(\Selector13~0_combout ),
	.cout());
defparam \Selector13~0 .lut_mask = 16'hE5E0;
defparam \Selector13~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_mem~19 (
	.dataa(csr_flash_cmd_addr_data_27),
	.datab(in_cmd_channel[1]),
	.datac(has_addr),
	.datad(in_cmd_channel[0]),
	.cin(gnd),
	.combout(\addr_mem~19_combout ),
	.cout());
defparam \addr_mem~19 .lut_mask = 16'h0080;
defparam \addr_mem~19 .sum_lutc_input = "datac";

dffeas \addr_mem[3][3] (
	.clk(clk_clk),
	.d(\addr_mem~19_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[3][3]~q ),
	.prn(vcc));
defparam \addr_mem[3][3] .is_wysiwyg = "true";
defparam \addr_mem[3][3] .power_up = "low";

cycloneive_lcell_comb \Selector13~1 (
	.dataa(\addr_mem[2][3]~q ),
	.datab(\addr_cnt[1]~q ),
	.datac(\Selector13~0_combout ),
	.datad(\addr_mem[3][3]~q ),
	.cin(gnd),
	.combout(\Selector13~1_combout ),
	.cout());
defparam \Selector13~1 .lut_mask = 16'hF838;
defparam \Selector13~1 .sum_lutc_input = "datac";

dffeas \header_information[3] (
	.clk(clk_clk),
	.d(in_cmd_data[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\header_information[3]~q ),
	.prn(vcc));
defparam \header_information[3] .is_wysiwyg = "true";
defparam \header_information[3] .power_up = "low";

cycloneive_lcell_comb \Selector13~2 (
	.dataa(\Selector13~1_combout ),
	.datab(\header_information[3]~q ),
	.datac(stateST_SEND_ADDR),
	.datad(\Selector9~0_combout ),
	.cin(gnd),
	.combout(\Selector13~2_combout ),
	.cout());
defparam \Selector13~2 .lut_mask = 16'h00AC;
defparam \Selector13~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_mem~20 (
	.dataa(csr_flash_cmd_addr_data_21),
	.datab(has_addr),
	.datac(mem_addr_reg_19),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\addr_mem~20_combout ),
	.cout());
defparam \addr_mem~20 .lut_mask = 16'h88F0;
defparam \addr_mem~20 .sum_lutc_input = "datac";

dffeas \addr_mem[2][5] (
	.clk(clk_clk),
	.d(\addr_mem~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[2][5]~q ),
	.prn(vcc));
defparam \addr_mem[2][5] .is_wysiwyg = "true";
defparam \addr_mem[2][5] .power_up = "low";

cycloneive_lcell_comb \addr_mem~21 (
	.dataa(csr_flash_cmd_addr_data_13),
	.datab(has_addr),
	.datac(mem_addr_reg_11),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\addr_mem~21_combout ),
	.cout());
defparam \addr_mem~21 .lut_mask = 16'h88F0;
defparam \addr_mem~21 .sum_lutc_input = "datac";

dffeas \addr_mem[1][5] (
	.clk(clk_clk),
	.d(\addr_mem~21_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[1][5]~q ),
	.prn(vcc));
defparam \addr_mem[1][5] .is_wysiwyg = "true";
defparam \addr_mem[1][5] .power_up = "low";

cycloneive_lcell_comb \addr_mem~22 (
	.dataa(csr_flash_cmd_addr_data_5),
	.datab(has_addr),
	.datac(mem_addr_reg_3),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\addr_mem~22_combout ),
	.cout());
defparam \addr_mem~22 .lut_mask = 16'h88F0;
defparam \addr_mem~22 .sum_lutc_input = "datac";

dffeas \addr_mem[0][5] (
	.clk(clk_clk),
	.d(\addr_mem~22_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[0][5]~q ),
	.prn(vcc));
defparam \addr_mem[0][5] .is_wysiwyg = "true";
defparam \addr_mem[0][5] .power_up = "low";

cycloneive_lcell_comb \Selector11~0 (
	.dataa(\addr_cnt[1]~q ),
	.datab(\addr_mem[1][5]~q ),
	.datac(\addr_cnt[0]~q ),
	.datad(\addr_mem[0][5]~q ),
	.cin(gnd),
	.combout(\Selector11~0_combout ),
	.cout());
defparam \Selector11~0 .lut_mask = 16'hE5E0;
defparam \Selector11~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_mem~23 (
	.dataa(csr_flash_cmd_addr_data_29),
	.datab(in_cmd_channel[1]),
	.datac(has_addr),
	.datad(in_cmd_channel[0]),
	.cin(gnd),
	.combout(\addr_mem~23_combout ),
	.cout());
defparam \addr_mem~23 .lut_mask = 16'h0080;
defparam \addr_mem~23 .sum_lutc_input = "datac";

dffeas \addr_mem[3][5] (
	.clk(clk_clk),
	.d(\addr_mem~23_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[3][5]~q ),
	.prn(vcc));
defparam \addr_mem[3][5] .is_wysiwyg = "true";
defparam \addr_mem[3][5] .power_up = "low";

cycloneive_lcell_comb \Selector11~1 (
	.dataa(\addr_mem[2][5]~q ),
	.datab(\addr_cnt[1]~q ),
	.datac(\Selector11~0_combout ),
	.datad(\addr_mem[3][5]~q ),
	.cin(gnd),
	.combout(\Selector11~1_combout ),
	.cout());
defparam \Selector11~1 .lut_mask = 16'hF838;
defparam \Selector11~1 .sum_lutc_input = "datac";

dffeas \header_information[5] (
	.clk(clk_clk),
	.d(in_cmd_data[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\header_information[5]~q ),
	.prn(vcc));
defparam \header_information[5] .is_wysiwyg = "true";
defparam \header_information[5] .power_up = "low";

cycloneive_lcell_comb \Selector11~2 (
	.dataa(\Selector11~1_combout ),
	.datab(\header_information[5]~q ),
	.datac(stateST_SEND_ADDR),
	.datad(\Selector9~0_combout ),
	.cin(gnd),
	.combout(\Selector11~2_combout ),
	.cout());
defparam \Selector11~2 .lut_mask = 16'h00AC;
defparam \Selector11~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_mem~24 (
	.dataa(csr_flash_cmd_addr_data_14),
	.datab(has_addr),
	.datac(mem_addr_reg_12),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\addr_mem~24_combout ),
	.cout());
defparam \addr_mem~24 .lut_mask = 16'h88F0;
defparam \addr_mem~24 .sum_lutc_input = "datac";

dffeas \addr_mem[1][6] (
	.clk(clk_clk),
	.d(\addr_mem~24_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[1][6]~q ),
	.prn(vcc));
defparam \addr_mem[1][6] .is_wysiwyg = "true";
defparam \addr_mem[1][6] .power_up = "low";

cycloneive_lcell_comb \addr_mem~25 (
	.dataa(csr_flash_cmd_addr_data_22),
	.datab(has_addr),
	.datac(mem_addr_reg_20),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\addr_mem~25_combout ),
	.cout());
defparam \addr_mem~25 .lut_mask = 16'h88F0;
defparam \addr_mem~25 .sum_lutc_input = "datac";

dffeas \addr_mem[2][6] (
	.clk(clk_clk),
	.d(\addr_mem~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[2][6]~q ),
	.prn(vcc));
defparam \addr_mem[2][6] .is_wysiwyg = "true";
defparam \addr_mem[2][6] .power_up = "low";

cycloneive_lcell_comb \addr_mem~26 (
	.dataa(csr_flash_cmd_addr_data_6),
	.datab(has_addr),
	.datac(mem_addr_reg_4),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\addr_mem~26_combout ),
	.cout());
defparam \addr_mem~26 .lut_mask = 16'h88F0;
defparam \addr_mem~26 .sum_lutc_input = "datac";

dffeas \addr_mem[0][6] (
	.clk(clk_clk),
	.d(\addr_mem~26_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[0][6]~q ),
	.prn(vcc));
defparam \addr_mem[0][6] .is_wysiwyg = "true";
defparam \addr_mem[0][6] .power_up = "low";

cycloneive_lcell_comb \Selector10~0 (
	.dataa(\addr_cnt[0]~q ),
	.datab(\addr_mem[2][6]~q ),
	.datac(\addr_cnt[1]~q ),
	.datad(\addr_mem[0][6]~q ),
	.cin(gnd),
	.combout(\Selector10~0_combout ),
	.cout());
defparam \Selector10~0 .lut_mask = 16'hE5E0;
defparam \Selector10~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_mem~27 (
	.dataa(csr_flash_cmd_addr_data_30),
	.datab(in_cmd_channel[1]),
	.datac(has_addr),
	.datad(in_cmd_channel[0]),
	.cin(gnd),
	.combout(\addr_mem~27_combout ),
	.cout());
defparam \addr_mem~27 .lut_mask = 16'h0080;
defparam \addr_mem~27 .sum_lutc_input = "datac";

dffeas \addr_mem[3][6] (
	.clk(clk_clk),
	.d(\addr_mem~27_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[3][6]~q ),
	.prn(vcc));
defparam \addr_mem[3][6] .is_wysiwyg = "true";
defparam \addr_mem[3][6] .power_up = "low";

cycloneive_lcell_comb \Selector10~1 (
	.dataa(\addr_mem[1][6]~q ),
	.datab(\addr_cnt[0]~q ),
	.datac(\Selector10~0_combout ),
	.datad(\addr_mem[3][6]~q ),
	.cin(gnd),
	.combout(\Selector10~1_combout ),
	.cout());
defparam \Selector10~1 .lut_mask = 16'hF838;
defparam \Selector10~1 .sum_lutc_input = "datac";

dffeas \header_information[6] (
	.clk(clk_clk),
	.d(in_cmd_data[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\header_information[6]~q ),
	.prn(vcc));
defparam \header_information[6] .is_wysiwyg = "true";
defparam \header_information[6] .power_up = "low";

cycloneive_lcell_comb \Selector10~2 (
	.dataa(\Selector10~1_combout ),
	.datab(stateST_SEND_OPCODE),
	.datac(\header_information[6]~q ),
	.datad(stateST_SEND_ADDR),
	.cin(gnd),
	.combout(\Selector10~2_combout ),
	.cout());
defparam \Selector10~2 .lut_mask = 16'hAAC0;
defparam \Selector10~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_mem~28 (
	.dataa(csr_flash_cmd_addr_data_23),
	.datab(in_cmd_channel[1]),
	.datac(has_addr),
	.datad(in_cmd_channel[0]),
	.cin(gnd),
	.combout(\addr_mem~28_combout ),
	.cout());
defparam \addr_mem~28 .lut_mask = 16'h0080;
defparam \addr_mem~28 .sum_lutc_input = "datac";

dffeas \addr_mem[2][7] (
	.clk(clk_clk),
	.d(\addr_mem~28_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[2][7]~q ),
	.prn(vcc));
defparam \addr_mem[2][7] .is_wysiwyg = "true";
defparam \addr_mem[2][7] .power_up = "low";

cycloneive_lcell_comb \addr_mem~29 (
	.dataa(csr_flash_cmd_addr_data_15),
	.datab(has_addr),
	.datac(mem_addr_reg_13),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\addr_mem~29_combout ),
	.cout());
defparam \addr_mem~29 .lut_mask = 16'h88F0;
defparam \addr_mem~29 .sum_lutc_input = "datac";

dffeas \addr_mem[1][7] (
	.clk(clk_clk),
	.d(\addr_mem~29_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[1][7]~q ),
	.prn(vcc));
defparam \addr_mem[1][7] .is_wysiwyg = "true";
defparam \addr_mem[1][7] .power_up = "low";

cycloneive_lcell_comb \addr_mem~30 (
	.dataa(csr_flash_cmd_addr_data_7),
	.datab(has_addr),
	.datac(mem_addr_reg_5),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\addr_mem~30_combout ),
	.cout());
defparam \addr_mem~30 .lut_mask = 16'h88F0;
defparam \addr_mem~30 .sum_lutc_input = "datac";

dffeas \addr_mem[0][7] (
	.clk(clk_clk),
	.d(\addr_mem~30_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[0][7]~q ),
	.prn(vcc));
defparam \addr_mem[0][7] .is_wysiwyg = "true";
defparam \addr_mem[0][7] .power_up = "low";

cycloneive_lcell_comb \Selector9~1 (
	.dataa(\addr_cnt[1]~q ),
	.datab(\addr_mem[1][7]~q ),
	.datac(\addr_cnt[0]~q ),
	.datad(\addr_mem[0][7]~q ),
	.cin(gnd),
	.combout(\Selector9~1_combout ),
	.cout());
defparam \Selector9~1 .lut_mask = 16'hE5E0;
defparam \Selector9~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \addr_mem~31 (
	.dataa(csr_flash_cmd_addr_data_31),
	.datab(in_cmd_channel[1]),
	.datac(has_addr),
	.datad(in_cmd_channel[0]),
	.cin(gnd),
	.combout(\addr_mem~31_combout ),
	.cout());
defparam \addr_mem~31 .lut_mask = 16'h0080;
defparam \addr_mem~31 .sum_lutc_input = "datac";

dffeas \addr_mem[3][7] (
	.clk(clk_clk),
	.d(\addr_mem~31_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\addr_mem[3][7]~q ),
	.prn(vcc));
defparam \addr_mem[3][7] .is_wysiwyg = "true";
defparam \addr_mem[3][7] .power_up = "low";

cycloneive_lcell_comb \Selector9~2 (
	.dataa(\addr_mem[2][7]~q ),
	.datab(\addr_cnt[1]~q ),
	.datac(\Selector9~1_combout ),
	.datad(\addr_mem[3][7]~q ),
	.cin(gnd),
	.combout(\Selector9~2_combout ),
	.cout());
defparam \Selector9~2 .lut_mask = 16'hF838;
defparam \Selector9~2 .sum_lutc_input = "datac";

dffeas \header_information[7] (
	.clk(clk_clk),
	.d(in_cmd_data[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\header_information[7]~q ),
	.prn(vcc));
defparam \header_information[7] .is_wysiwyg = "true";
defparam \header_information[7] .power_up = "low";

cycloneive_lcell_comb \Selector9~3 (
	.dataa(\Selector9~2_combout ),
	.datab(\header_information[7]~q ),
	.datac(stateST_SEND_ADDR),
	.datad(\Selector9~0_combout ),
	.cin(gnd),
	.combout(\Selector9~3_combout ),
	.cout());
defparam \Selector9~3 .lut_mask = 16'h00AC;
defparam \Selector9~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector3~5 (
	.dataa(stateST_SEND_OPCODE),
	.datab(gnd),
	.datac(gnd),
	.datad(\header_information[8]~q ),
	.cin(gnd),
	.combout(\Selector3~5_combout ),
	.cout());
defparam \Selector3~5 .lut_mask = 16'h00AA;
defparam \Selector3~5 .sum_lutc_input = "datac";

endmodule

module flashLoader_data_adapter_32_8 (
	reset,
	state_register_1,
	state_register_0,
	out_valid1,
	a_valid1,
	stateST_SEND_DATA,
	WideOr0,
	WideOr01,
	in_valid,
	out_data_0,
	out_data_4,
	out_data_2,
	out_data_1,
	out_data_3,
	out_data_5,
	out_data_6,
	out_data_7,
	in_data,
	clk)/* synthesis synthesis_greybox=0 */;
input 	reset;
output 	state_register_1;
output 	state_register_0;
output 	out_valid1;
output 	a_valid1;
input 	stateST_SEND_DATA;
input 	WideOr0;
input 	WideOr01;
input 	in_valid;
output 	out_data_0;
output 	out_data_4;
output 	out_data_2;
output 	out_data_1;
output 	out_data_3;
output 	out_data_5;
output 	out_data_6;
output 	out_data_7;
input 	[31:0] in_data;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always4~0_combout ;
wire \Mux9~0_combout ;
wire \state_register[0]~0_combout ;
wire \in_ready~0_combout ;
wire \in_ready~1_combout ;
wire \a_data1[0]~q ;
wire \a_data2[0]~q ;
wire \a_data0[0]~q ;
wire \Mux7~0_combout ;
wire \a_data3[0]~q ;
wire \Mux7~1_combout ;
wire \a_data1[4]~q ;
wire \a_data2[4]~q ;
wire \a_data0[4]~q ;
wire \Mux3~0_combout ;
wire \a_data3[4]~q ;
wire \Mux3~1_combout ;
wire \a_data1[2]~q ;
wire \a_data2[2]~q ;
wire \a_data0[2]~q ;
wire \Mux5~0_combout ;
wire \a_data3[2]~q ;
wire \Mux5~1_combout ;
wire \a_data2[1]~q ;
wire \a_data1[1]~q ;
wire \a_data0[1]~q ;
wire \Mux6~0_combout ;
wire \a_data3[1]~q ;
wire \Mux6~1_combout ;
wire \a_data2[3]~q ;
wire \a_data1[3]~q ;
wire \a_data0[3]~q ;
wire \Mux4~0_combout ;
wire \a_data3[3]~q ;
wire \Mux4~1_combout ;
wire \a_data2[5]~q ;
wire \a_data1[5]~q ;
wire \a_data0[5]~q ;
wire \Mux2~0_combout ;
wire \a_data3[5]~q ;
wire \Mux2~1_combout ;
wire \a_data1[6]~q ;
wire \a_data2[6]~q ;
wire \a_data0[6]~q ;
wire \Mux1~0_combout ;
wire \a_data3[6]~q ;
wire \Mux1~1_combout ;
wire \a_data2[7]~q ;
wire \a_data1[7]~q ;
wire \a_data0[7]~q ;
wire \Mux0~0_combout ;
wire \a_data3[7]~q ;
wire \Mux0~1_combout ;


dffeas \state_register[1] (
	.clk(clk),
	.d(\Mux9~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(state_register_1),
	.prn(vcc));
defparam \state_register[1] .is_wysiwyg = "true";
defparam \state_register[1] .power_up = "low";

dffeas \state_register[0] (
	.clk(clk),
	.d(\state_register[0]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(state_register_0),
	.prn(vcc));
defparam \state_register[0] .is_wysiwyg = "true";
defparam \state_register[0] .power_up = "low";

dffeas out_valid(
	.clk(clk),
	.d(a_valid1),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(out_valid1),
	.prn(vcc));
defparam out_valid.is_wysiwyg = "true";
defparam out_valid.power_up = "low";

dffeas a_valid(
	.clk(clk),
	.d(in_valid),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(a_valid1),
	.prn(vcc));
defparam a_valid.is_wysiwyg = "true";
defparam a_valid.power_up = "low";

dffeas \out_data[0] (
	.clk(clk),
	.d(\Mux7~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(out_data_0),
	.prn(vcc));
defparam \out_data[0] .is_wysiwyg = "true";
defparam \out_data[0] .power_up = "low";

dffeas \out_data[4] (
	.clk(clk),
	.d(\Mux3~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(out_data_4),
	.prn(vcc));
defparam \out_data[4] .is_wysiwyg = "true";
defparam \out_data[4] .power_up = "low";

dffeas \out_data[2] (
	.clk(clk),
	.d(\Mux5~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(out_data_2),
	.prn(vcc));
defparam \out_data[2] .is_wysiwyg = "true";
defparam \out_data[2] .power_up = "low";

dffeas \out_data[1] (
	.clk(clk),
	.d(\Mux6~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(out_data_1),
	.prn(vcc));
defparam \out_data[1] .is_wysiwyg = "true";
defparam \out_data[1] .power_up = "low";

dffeas \out_data[3] (
	.clk(clk),
	.d(\Mux4~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(out_data_3),
	.prn(vcc));
defparam \out_data[3] .is_wysiwyg = "true";
defparam \out_data[3] .power_up = "low";

dffeas \out_data[5] (
	.clk(clk),
	.d(\Mux2~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(out_data_5),
	.prn(vcc));
defparam \out_data[5] .is_wysiwyg = "true";
defparam \out_data[5] .power_up = "low";

dffeas \out_data[6] (
	.clk(clk),
	.d(\Mux1~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(out_data_6),
	.prn(vcc));
defparam \out_data[6] .is_wysiwyg = "true";
defparam \out_data[6] .power_up = "low";

dffeas \out_data[7] (
	.clk(clk),
	.d(\Mux0~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~0_combout ),
	.q(out_data_7),
	.prn(vcc));
defparam \out_data[7] .is_wysiwyg = "true";
defparam \out_data[7] .power_up = "low";

cycloneive_lcell_comb \always4~0 (
	.dataa(stateST_SEND_DATA),
	.datab(WideOr01),
	.datac(WideOr0),
	.datad(out_valid1),
	.cin(gnd),
	.combout(\always4~0_combout ),
	.cout());
defparam \always4~0 .lut_mask = 16'hA8FF;
defparam \always4~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux9~0 (
	.dataa(state_register_1),
	.datab(state_register_0),
	.datac(a_valid1),
	.datad(\always4~0_combout ),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
defparam \Mux9~0 .lut_mask = 16'h6AAA;
defparam \Mux9~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \state_register[0]~0 (
	.dataa(gnd),
	.datab(state_register_0),
	.datac(a_valid1),
	.datad(\always4~0_combout ),
	.cin(gnd),
	.combout(\state_register[0]~0_combout ),
	.cout());
defparam \state_register[0]~0 .lut_mask = 16'h3CCC;
defparam \state_register[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \in_ready~0 (
	.dataa(stateST_SEND_DATA),
	.datab(out_valid1),
	.datac(WideOr01),
	.datad(WideOr0),
	.cin(gnd),
	.combout(\in_ready~0_combout ),
	.cout());
defparam \in_ready~0 .lut_mask = 16'h444C;
defparam \in_ready~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \in_ready~1 (
	.dataa(state_register_1),
	.datab(state_register_0),
	.datac(a_valid1),
	.datad(\in_ready~0_combout ),
	.cin(gnd),
	.combout(\in_ready~1_combout ),
	.cout());
defparam \in_ready~1 .lut_mask = 16'h0F8F;
defparam \in_ready~1 .sum_lutc_input = "datac";

dffeas \a_data1[0] (
	.clk(clk),
	.d(in_data[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data1[0]~q ),
	.prn(vcc));
defparam \a_data1[0] .is_wysiwyg = "true";
defparam \a_data1[0] .power_up = "low";

dffeas \a_data2[0] (
	.clk(clk),
	.d(in_data[16]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data2[0]~q ),
	.prn(vcc));
defparam \a_data2[0] .is_wysiwyg = "true";
defparam \a_data2[0] .power_up = "low";

dffeas \a_data0[0] (
	.clk(clk),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data0[0]~q ),
	.prn(vcc));
defparam \a_data0[0] .is_wysiwyg = "true";
defparam \a_data0[0] .power_up = "low";

cycloneive_lcell_comb \Mux7~0 (
	.dataa(state_register_0),
	.datab(\a_data2[0]~q ),
	.datac(state_register_1),
	.datad(\a_data0[0]~q ),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
defparam \Mux7~0 .lut_mask = 16'hE5E0;
defparam \Mux7~0 .sum_lutc_input = "datac";

dffeas \a_data3[0] (
	.clk(clk),
	.d(in_data[24]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data3[0]~q ),
	.prn(vcc));
defparam \a_data3[0] .is_wysiwyg = "true";
defparam \a_data3[0] .power_up = "low";

cycloneive_lcell_comb \Mux7~1 (
	.dataa(\a_data1[0]~q ),
	.datab(state_register_0),
	.datac(\Mux7~0_combout ),
	.datad(\a_data3[0]~q ),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
defparam \Mux7~1 .lut_mask = 16'hF838;
defparam \Mux7~1 .sum_lutc_input = "datac";

dffeas \a_data1[4] (
	.clk(clk),
	.d(in_data[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data1[4]~q ),
	.prn(vcc));
defparam \a_data1[4] .is_wysiwyg = "true";
defparam \a_data1[4] .power_up = "low";

dffeas \a_data2[4] (
	.clk(clk),
	.d(in_data[20]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data2[4]~q ),
	.prn(vcc));
defparam \a_data2[4] .is_wysiwyg = "true";
defparam \a_data2[4] .power_up = "low";

dffeas \a_data0[4] (
	.clk(clk),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data0[4]~q ),
	.prn(vcc));
defparam \a_data0[4] .is_wysiwyg = "true";
defparam \a_data0[4] .power_up = "low";

cycloneive_lcell_comb \Mux3~0 (
	.dataa(state_register_0),
	.datab(\a_data2[4]~q ),
	.datac(state_register_1),
	.datad(\a_data0[4]~q ),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'hE5E0;
defparam \Mux3~0 .sum_lutc_input = "datac";

dffeas \a_data3[4] (
	.clk(clk),
	.d(in_data[28]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data3[4]~q ),
	.prn(vcc));
defparam \a_data3[4] .is_wysiwyg = "true";
defparam \a_data3[4] .power_up = "low";

cycloneive_lcell_comb \Mux3~1 (
	.dataa(\a_data1[4]~q ),
	.datab(state_register_0),
	.datac(\Mux3~0_combout ),
	.datad(\a_data3[4]~q ),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
defparam \Mux3~1 .lut_mask = 16'hF838;
defparam \Mux3~1 .sum_lutc_input = "datac";

dffeas \a_data1[2] (
	.clk(clk),
	.d(in_data[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data1[2]~q ),
	.prn(vcc));
defparam \a_data1[2] .is_wysiwyg = "true";
defparam \a_data1[2] .power_up = "low";

dffeas \a_data2[2] (
	.clk(clk),
	.d(in_data[18]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data2[2]~q ),
	.prn(vcc));
defparam \a_data2[2] .is_wysiwyg = "true";
defparam \a_data2[2] .power_up = "low";

dffeas \a_data0[2] (
	.clk(clk),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data0[2]~q ),
	.prn(vcc));
defparam \a_data0[2] .is_wysiwyg = "true";
defparam \a_data0[2] .power_up = "low";

cycloneive_lcell_comb \Mux5~0 (
	.dataa(state_register_0),
	.datab(\a_data2[2]~q ),
	.datac(state_register_1),
	.datad(\a_data0[2]~q ),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
defparam \Mux5~0 .lut_mask = 16'hE5E0;
defparam \Mux5~0 .sum_lutc_input = "datac";

dffeas \a_data3[2] (
	.clk(clk),
	.d(in_data[26]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data3[2]~q ),
	.prn(vcc));
defparam \a_data3[2] .is_wysiwyg = "true";
defparam \a_data3[2] .power_up = "low";

cycloneive_lcell_comb \Mux5~1 (
	.dataa(\a_data1[2]~q ),
	.datab(state_register_0),
	.datac(\Mux5~0_combout ),
	.datad(\a_data3[2]~q ),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
defparam \Mux5~1 .lut_mask = 16'hF838;
defparam \Mux5~1 .sum_lutc_input = "datac";

dffeas \a_data2[1] (
	.clk(clk),
	.d(in_data[17]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data2[1]~q ),
	.prn(vcc));
defparam \a_data2[1] .is_wysiwyg = "true";
defparam \a_data2[1] .power_up = "low";

dffeas \a_data1[1] (
	.clk(clk),
	.d(in_data[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data1[1]~q ),
	.prn(vcc));
defparam \a_data1[1] .is_wysiwyg = "true";
defparam \a_data1[1] .power_up = "low";

dffeas \a_data0[1] (
	.clk(clk),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data0[1]~q ),
	.prn(vcc));
defparam \a_data0[1] .is_wysiwyg = "true";
defparam \a_data0[1] .power_up = "low";

cycloneive_lcell_comb \Mux6~0 (
	.dataa(state_register_1),
	.datab(\a_data1[1]~q ),
	.datac(state_register_0),
	.datad(\a_data0[1]~q ),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
defparam \Mux6~0 .lut_mask = 16'hE5E0;
defparam \Mux6~0 .sum_lutc_input = "datac";

dffeas \a_data3[1] (
	.clk(clk),
	.d(in_data[25]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data3[1]~q ),
	.prn(vcc));
defparam \a_data3[1] .is_wysiwyg = "true";
defparam \a_data3[1] .power_up = "low";

cycloneive_lcell_comb \Mux6~1 (
	.dataa(\a_data2[1]~q ),
	.datab(state_register_1),
	.datac(\Mux6~0_combout ),
	.datad(\a_data3[1]~q ),
	.cin(gnd),
	.combout(\Mux6~1_combout ),
	.cout());
defparam \Mux6~1 .lut_mask = 16'hF838;
defparam \Mux6~1 .sum_lutc_input = "datac";

dffeas \a_data2[3] (
	.clk(clk),
	.d(in_data[19]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data2[3]~q ),
	.prn(vcc));
defparam \a_data2[3] .is_wysiwyg = "true";
defparam \a_data2[3] .power_up = "low";

dffeas \a_data1[3] (
	.clk(clk),
	.d(in_data[11]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data1[3]~q ),
	.prn(vcc));
defparam \a_data1[3] .is_wysiwyg = "true";
defparam \a_data1[3] .power_up = "low";

dffeas \a_data0[3] (
	.clk(clk),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data0[3]~q ),
	.prn(vcc));
defparam \a_data0[3] .is_wysiwyg = "true";
defparam \a_data0[3] .power_up = "low";

cycloneive_lcell_comb \Mux4~0 (
	.dataa(state_register_1),
	.datab(\a_data1[3]~q ),
	.datac(state_register_0),
	.datad(\a_data0[3]~q ),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
defparam \Mux4~0 .lut_mask = 16'hE5E0;
defparam \Mux4~0 .sum_lutc_input = "datac";

dffeas \a_data3[3] (
	.clk(clk),
	.d(in_data[27]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data3[3]~q ),
	.prn(vcc));
defparam \a_data3[3] .is_wysiwyg = "true";
defparam \a_data3[3] .power_up = "low";

cycloneive_lcell_comb \Mux4~1 (
	.dataa(\a_data2[3]~q ),
	.datab(state_register_1),
	.datac(\Mux4~0_combout ),
	.datad(\a_data3[3]~q ),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
defparam \Mux4~1 .lut_mask = 16'hF838;
defparam \Mux4~1 .sum_lutc_input = "datac";

dffeas \a_data2[5] (
	.clk(clk),
	.d(in_data[21]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data2[5]~q ),
	.prn(vcc));
defparam \a_data2[5] .is_wysiwyg = "true";
defparam \a_data2[5] .power_up = "low";

dffeas \a_data1[5] (
	.clk(clk),
	.d(in_data[13]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data1[5]~q ),
	.prn(vcc));
defparam \a_data1[5] .is_wysiwyg = "true";
defparam \a_data1[5] .power_up = "low";

dffeas \a_data0[5] (
	.clk(clk),
	.d(in_data[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data0[5]~q ),
	.prn(vcc));
defparam \a_data0[5] .is_wysiwyg = "true";
defparam \a_data0[5] .power_up = "low";

cycloneive_lcell_comb \Mux2~0 (
	.dataa(state_register_1),
	.datab(\a_data1[5]~q ),
	.datac(state_register_0),
	.datad(\a_data0[5]~q ),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
defparam \Mux2~0 .lut_mask = 16'hE5E0;
defparam \Mux2~0 .sum_lutc_input = "datac";

dffeas \a_data3[5] (
	.clk(clk),
	.d(in_data[29]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data3[5]~q ),
	.prn(vcc));
defparam \a_data3[5] .is_wysiwyg = "true";
defparam \a_data3[5] .power_up = "low";

cycloneive_lcell_comb \Mux2~1 (
	.dataa(\a_data2[5]~q ),
	.datab(state_register_1),
	.datac(\Mux2~0_combout ),
	.datad(\a_data3[5]~q ),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
defparam \Mux2~1 .lut_mask = 16'hF838;
defparam \Mux2~1 .sum_lutc_input = "datac";

dffeas \a_data1[6] (
	.clk(clk),
	.d(in_data[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data1[6]~q ),
	.prn(vcc));
defparam \a_data1[6] .is_wysiwyg = "true";
defparam \a_data1[6] .power_up = "low";

dffeas \a_data2[6] (
	.clk(clk),
	.d(in_data[22]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data2[6]~q ),
	.prn(vcc));
defparam \a_data2[6] .is_wysiwyg = "true";
defparam \a_data2[6] .power_up = "low";

dffeas \a_data0[6] (
	.clk(clk),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data0[6]~q ),
	.prn(vcc));
defparam \a_data0[6] .is_wysiwyg = "true";
defparam \a_data0[6] .power_up = "low";

cycloneive_lcell_comb \Mux1~0 (
	.dataa(state_register_0),
	.datab(\a_data2[6]~q ),
	.datac(state_register_1),
	.datad(\a_data0[6]~q ),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'hE5E0;
defparam \Mux1~0 .sum_lutc_input = "datac";

dffeas \a_data3[6] (
	.clk(clk),
	.d(in_data[30]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data3[6]~q ),
	.prn(vcc));
defparam \a_data3[6] .is_wysiwyg = "true";
defparam \a_data3[6] .power_up = "low";

cycloneive_lcell_comb \Mux1~1 (
	.dataa(\a_data1[6]~q ),
	.datab(state_register_0),
	.datac(\Mux1~0_combout ),
	.datad(\a_data3[6]~q ),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
defparam \Mux1~1 .lut_mask = 16'hF838;
defparam \Mux1~1 .sum_lutc_input = "datac";

dffeas \a_data2[7] (
	.clk(clk),
	.d(in_data[23]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data2[7]~q ),
	.prn(vcc));
defparam \a_data2[7] .is_wysiwyg = "true";
defparam \a_data2[7] .power_up = "low";

dffeas \a_data1[7] (
	.clk(clk),
	.d(in_data[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data1[7]~q ),
	.prn(vcc));
defparam \a_data1[7] .is_wysiwyg = "true";
defparam \a_data1[7] .power_up = "low";

dffeas \a_data0[7] (
	.clk(clk),
	.d(in_data[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data0[7]~q ),
	.prn(vcc));
defparam \a_data0[7] .is_wysiwyg = "true";
defparam \a_data0[7] .power_up = "low";

cycloneive_lcell_comb \Mux0~0 (
	.dataa(state_register_1),
	.datab(\a_data1[7]~q ),
	.datac(state_register_0),
	.datad(\a_data0[7]~q ),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hE5E0;
defparam \Mux0~0 .sum_lutc_input = "datac";

dffeas \a_data3[7] (
	.clk(clk),
	.d(in_data[31]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~1_combout ),
	.q(\a_data3[7]~q ),
	.prn(vcc));
defparam \a_data3[7] .is_wysiwyg = "true";
defparam \a_data3[7] .power_up = "low";

cycloneive_lcell_comb \Mux0~1 (
	.dataa(\a_data2[7]~q ),
	.datab(state_register_1),
	.datac(\Mux0~0_combout ),
	.datad(\a_data3[7]~q ),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hF838;
defparam \Mux0~1 .sum_lutc_input = "datac";

endmodule

module flashLoader_data_adapter_8_32 (
	out_valid1,
	out_endofpacket1,
	in_cmd_channel_reg_1,
	stateST_WAIT_RSP,
	out_data_0,
	out_data_1,
	out_data_2,
	out_data_3,
	out_data_4,
	out_data_5,
	out_data_6,
	out_data_7,
	out_data_8,
	out_data_9,
	out_data_10,
	out_data_11,
	out_data_12,
	out_data_13,
	out_data_14,
	out_data_15,
	out_data_16,
	out_data_17,
	out_data_18,
	out_data_19,
	out_data_20,
	out_data_21,
	out_data_22,
	out_data_23,
	out_data_24,
	out_data_25,
	out_data_26,
	out_data_27,
	out_data_28,
	out_data_29,
	out_data_30,
	out_data_31,
	in_cmd_channel_reg_0,
	a_valid1,
	a_ready1,
	reset,
	in_valid,
	in_ready1,
	in_endofpacket,
	in_data,
	clk)/* synthesis synthesis_greybox=0 */;
output 	out_valid1;
output 	out_endofpacket1;
input 	in_cmd_channel_reg_1;
input 	stateST_WAIT_RSP;
output 	out_data_0;
output 	out_data_1;
output 	out_data_2;
output 	out_data_3;
output 	out_data_4;
output 	out_data_5;
output 	out_data_6;
output 	out_data_7;
output 	out_data_8;
output 	out_data_9;
output 	out_data_10;
output 	out_data_11;
output 	out_data_12;
output 	out_data_13;
output 	out_data_14;
output 	out_data_15;
output 	out_data_16;
output 	out_data_17;
output 	out_data_18;
output 	out_data_19;
output 	out_data_20;
output 	out_data_21;
output 	out_data_22;
output 	out_data_23;
output 	out_data_24;
output 	out_data_25;
output 	out_data_26;
output 	out_data_27;
output 	out_data_28;
output 	out_data_29;
output 	out_data_30;
output 	out_data_31;
input 	in_cmd_channel_reg_0;
output 	a_valid1;
output 	a_ready1;
input 	reset;
input 	in_valid;
output 	in_ready1;
input 	in_endofpacket;
input 	[7:0] in_data;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a_endofpacket~q ;
wire \Mux17~0_combout ;
wire \state_register[0]~q ;
wire \state_d1[0]~q ;
wire \in_ready_d1~q ;
wire \state[0]~0_combout ;
wire \new_state~0_combout ;
wire \Mux16~0_combout ;
wire \state_register[1]~q ;
wire \state_d1[1]~q ;
wire \state[1]~1_combout ;
wire \out_valid~0_combout ;
wire \out_valid~1_combout ;
wire \a_data0[0]~q ;
wire \data0_register[0]~0_combout ;
wire \data0_register[0]~q ;
wire \b_data[0]~0_combout ;
wire \a_data0[1]~q ;
wire \data0_register[1]~q ;
wire \b_data[1]~1_combout ;
wire \a_data0[2]~q ;
wire \data0_register[2]~q ;
wire \b_data[2]~2_combout ;
wire \a_data0[3]~q ;
wire \data0_register[3]~q ;
wire \b_data[3]~3_combout ;
wire \a_data0[4]~q ;
wire \data0_register[4]~q ;
wire \b_data[4]~4_combout ;
wire \a_data0[5]~q ;
wire \data0_register[5]~q ;
wire \b_data[5]~5_combout ;
wire \a_data0[6]~q ;
wire \data0_register[6]~q ;
wire \b_data[6]~6_combout ;
wire \a_data0[7]~q ;
wire \data0_register[7]~q ;
wire \b_data[7]~7_combout ;
wire \data1_register[0]~0_combout ;
wire \data1_register[0]~q ;
wire \Mux15~0_combout ;
wire \data1_register[1]~q ;
wire \Mux14~0_combout ;
wire \data1_register[2]~q ;
wire \Mux13~0_combout ;
wire \data1_register[3]~q ;
wire \Mux12~0_combout ;
wire \data1_register[4]~q ;
wire \Mux11~0_combout ;
wire \data1_register[5]~q ;
wire \Mux10~0_combout ;
wire \data1_register[6]~q ;
wire \Mux9~0_combout ;
wire \data1_register[7]~q ;
wire \Mux8~0_combout ;
wire \mem_write2~0_combout ;
wire \data2_register[0]~q ;
wire \Mux7~0_combout ;
wire \data2_register[1]~q ;
wire \Mux6~0_combout ;
wire \data2_register[2]~q ;
wire \Mux5~0_combout ;
wire \data2_register[3]~q ;
wire \Mux4~0_combout ;
wire \data2_register[4]~q ;
wire \Mux3~0_combout ;
wire \data2_register[5]~q ;
wire \Mux2~0_combout ;
wire \data2_register[6]~q ;
wire \Mux1~0_combout ;
wire \data2_register[7]~q ;
wire \Mux0~0_combout ;
wire \b_data[24]~8_combout ;
wire \b_data[25]~9_combout ;
wire \b_data[26]~10_combout ;
wire \b_data[27]~11_combout ;
wire \b_data[28]~12_combout ;
wire \b_data[29]~13_combout ;
wire \b_data[30]~14_combout ;
wire \b_data[31]~15_combout ;


dffeas out_valid(
	.clk(clk),
	.d(\out_valid~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_valid1),
	.prn(vcc));
defparam out_valid.is_wysiwyg = "true";
defparam out_valid.power_up = "low";

dffeas out_endofpacket(
	.clk(clk),
	.d(\a_endofpacket~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_endofpacket1),
	.prn(vcc));
defparam out_endofpacket.is_wysiwyg = "true";
defparam out_endofpacket.power_up = "low";

dffeas \out_data[0] (
	.clk(clk),
	.d(\b_data[0]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_0),
	.prn(vcc));
defparam \out_data[0] .is_wysiwyg = "true";
defparam \out_data[0] .power_up = "low";

dffeas \out_data[1] (
	.clk(clk),
	.d(\b_data[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_1),
	.prn(vcc));
defparam \out_data[1] .is_wysiwyg = "true";
defparam \out_data[1] .power_up = "low";

dffeas \out_data[2] (
	.clk(clk),
	.d(\b_data[2]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_2),
	.prn(vcc));
defparam \out_data[2] .is_wysiwyg = "true";
defparam \out_data[2] .power_up = "low";

dffeas \out_data[3] (
	.clk(clk),
	.d(\b_data[3]~3_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_3),
	.prn(vcc));
defparam \out_data[3] .is_wysiwyg = "true";
defparam \out_data[3] .power_up = "low";

dffeas \out_data[4] (
	.clk(clk),
	.d(\b_data[4]~4_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_4),
	.prn(vcc));
defparam \out_data[4] .is_wysiwyg = "true";
defparam \out_data[4] .power_up = "low";

dffeas \out_data[5] (
	.clk(clk),
	.d(\b_data[5]~5_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_5),
	.prn(vcc));
defparam \out_data[5] .is_wysiwyg = "true";
defparam \out_data[5] .power_up = "low";

dffeas \out_data[6] (
	.clk(clk),
	.d(\b_data[6]~6_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_6),
	.prn(vcc));
defparam \out_data[6] .is_wysiwyg = "true";
defparam \out_data[6] .power_up = "low";

dffeas \out_data[7] (
	.clk(clk),
	.d(\b_data[7]~7_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_7),
	.prn(vcc));
defparam \out_data[7] .is_wysiwyg = "true";
defparam \out_data[7] .power_up = "low";

dffeas \out_data[8] (
	.clk(clk),
	.d(\Mux15~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_8),
	.prn(vcc));
defparam \out_data[8] .is_wysiwyg = "true";
defparam \out_data[8] .power_up = "low";

dffeas \out_data[9] (
	.clk(clk),
	.d(\Mux14~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_9),
	.prn(vcc));
defparam \out_data[9] .is_wysiwyg = "true";
defparam \out_data[9] .power_up = "low";

dffeas \out_data[10] (
	.clk(clk),
	.d(\Mux13~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_10),
	.prn(vcc));
defparam \out_data[10] .is_wysiwyg = "true";
defparam \out_data[10] .power_up = "low";

dffeas \out_data[11] (
	.clk(clk),
	.d(\Mux12~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_11),
	.prn(vcc));
defparam \out_data[11] .is_wysiwyg = "true";
defparam \out_data[11] .power_up = "low";

dffeas \out_data[12] (
	.clk(clk),
	.d(\Mux11~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_12),
	.prn(vcc));
defparam \out_data[12] .is_wysiwyg = "true";
defparam \out_data[12] .power_up = "low";

dffeas \out_data[13] (
	.clk(clk),
	.d(\Mux10~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_13),
	.prn(vcc));
defparam \out_data[13] .is_wysiwyg = "true";
defparam \out_data[13] .power_up = "low";

dffeas \out_data[14] (
	.clk(clk),
	.d(\Mux9~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_14),
	.prn(vcc));
defparam \out_data[14] .is_wysiwyg = "true";
defparam \out_data[14] .power_up = "low";

dffeas \out_data[15] (
	.clk(clk),
	.d(\Mux8~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_15),
	.prn(vcc));
defparam \out_data[15] .is_wysiwyg = "true";
defparam \out_data[15] .power_up = "low";

dffeas \out_data[16] (
	.clk(clk),
	.d(\Mux7~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_16),
	.prn(vcc));
defparam \out_data[16] .is_wysiwyg = "true";
defparam \out_data[16] .power_up = "low";

dffeas \out_data[17] (
	.clk(clk),
	.d(\Mux6~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_17),
	.prn(vcc));
defparam \out_data[17] .is_wysiwyg = "true";
defparam \out_data[17] .power_up = "low";

dffeas \out_data[18] (
	.clk(clk),
	.d(\Mux5~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_18),
	.prn(vcc));
defparam \out_data[18] .is_wysiwyg = "true";
defparam \out_data[18] .power_up = "low";

dffeas \out_data[19] (
	.clk(clk),
	.d(\Mux4~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_19),
	.prn(vcc));
defparam \out_data[19] .is_wysiwyg = "true";
defparam \out_data[19] .power_up = "low";

dffeas \out_data[20] (
	.clk(clk),
	.d(\Mux3~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_20),
	.prn(vcc));
defparam \out_data[20] .is_wysiwyg = "true";
defparam \out_data[20] .power_up = "low";

dffeas \out_data[21] (
	.clk(clk),
	.d(\Mux2~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_21),
	.prn(vcc));
defparam \out_data[21] .is_wysiwyg = "true";
defparam \out_data[21] .power_up = "low";

dffeas \out_data[22] (
	.clk(clk),
	.d(\Mux1~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_22),
	.prn(vcc));
defparam \out_data[22] .is_wysiwyg = "true";
defparam \out_data[22] .power_up = "low";

dffeas \out_data[23] (
	.clk(clk),
	.d(\Mux0~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_23),
	.prn(vcc));
defparam \out_data[23] .is_wysiwyg = "true";
defparam \out_data[23] .power_up = "low";

dffeas \out_data[24] (
	.clk(clk),
	.d(\b_data[24]~8_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_24),
	.prn(vcc));
defparam \out_data[24] .is_wysiwyg = "true";
defparam \out_data[24] .power_up = "low";

dffeas \out_data[25] (
	.clk(clk),
	.d(\b_data[25]~9_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_25),
	.prn(vcc));
defparam \out_data[25] .is_wysiwyg = "true";
defparam \out_data[25] .power_up = "low";

dffeas \out_data[26] (
	.clk(clk),
	.d(\b_data[26]~10_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_26),
	.prn(vcc));
defparam \out_data[26] .is_wysiwyg = "true";
defparam \out_data[26] .power_up = "low";

dffeas \out_data[27] (
	.clk(clk),
	.d(\b_data[27]~11_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_27),
	.prn(vcc));
defparam \out_data[27] .is_wysiwyg = "true";
defparam \out_data[27] .power_up = "low";

dffeas \out_data[28] (
	.clk(clk),
	.d(\b_data[28]~12_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_28),
	.prn(vcc));
defparam \out_data[28] .is_wysiwyg = "true";
defparam \out_data[28] .power_up = "low";

dffeas \out_data[29] (
	.clk(clk),
	.d(\b_data[29]~13_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_29),
	.prn(vcc));
defparam \out_data[29] .is_wysiwyg = "true";
defparam \out_data[29] .power_up = "low";

dffeas \out_data[30] (
	.clk(clk),
	.d(\b_data[30]~14_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_30),
	.prn(vcc));
defparam \out_data[30] .is_wysiwyg = "true";
defparam \out_data[30] .power_up = "low";

dffeas \out_data[31] (
	.clk(clk),
	.d(\b_data[31]~15_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(a_ready1),
	.q(out_data_31),
	.prn(vcc));
defparam \out_data[31] .is_wysiwyg = "true";
defparam \out_data[31] .power_up = "low";

dffeas a_valid(
	.clk(clk),
	.d(in_valid),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(a_valid1),
	.prn(vcc));
defparam a_valid.is_wysiwyg = "true";
defparam a_valid.power_up = "low";

cycloneive_lcell_comb a_ready(
	.dataa(in_cmd_channel_reg_0),
	.datab(in_cmd_channel_reg_1),
	.datac(stateST_WAIT_RSP),
	.datad(out_valid1),
	.cin(gnd),
	.combout(a_ready1),
	.cout());
defparam a_ready.lut_mask = 16'hEAFF;
defparam a_ready.sum_lutc_input = "datac";

cycloneive_lcell_comb in_ready(
	.dataa(a_ready1),
	.datab(gnd),
	.datac(gnd),
	.datad(a_valid1),
	.cin(gnd),
	.combout(in_ready1),
	.cout());
defparam in_ready.lut_mask = 16'hAAFF;
defparam in_ready.sum_lutc_input = "datac";

dffeas a_endofpacket(
	.clk(clk),
	.d(in_endofpacket),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_endofpacket~q ),
	.prn(vcc));
defparam a_endofpacket.is_wysiwyg = "true";
defparam a_endofpacket.power_up = "low";

cycloneive_lcell_comb \Mux17~0 (
	.dataa(a_ready1),
	.datab(a_valid1),
	.datac(\a_endofpacket~q ),
	.datad(\state[0]~0_combout ),
	.cin(gnd),
	.combout(\Mux17~0_combout ),
	.cout());
defparam \Mux17~0 .lut_mask = 16'h7708;
defparam \Mux17~0 .sum_lutc_input = "datac";

dffeas \state_register[0] (
	.clk(clk),
	.d(\Mux17~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state_register[0]~q ),
	.prn(vcc));
defparam \state_register[0] .is_wysiwyg = "true";
defparam \state_register[0] .power_up = "low";

dffeas \state_d1[0] (
	.clk(clk),
	.d(\state[0]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state_d1[0]~q ),
	.prn(vcc));
defparam \state_d1[0] .is_wysiwyg = "true";
defparam \state_d1[0] .power_up = "low";

dffeas in_ready_d1(
	.clk(clk),
	.d(in_ready1),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\in_ready_d1~q ),
	.prn(vcc));
defparam in_ready_d1.is_wysiwyg = "true";
defparam in_ready_d1.power_up = "low";

cycloneive_lcell_comb \state[0]~0 (
	.dataa(\state_register[0]~q ),
	.datab(\state_d1[0]~q ),
	.datac(gnd),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\state[0]~0_combout ),
	.cout());
defparam \state[0]~0 .lut_mask = 16'hAACC;
defparam \state[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \new_state~0 (
	.dataa(a_ready1),
	.datab(a_valid1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\new_state~0_combout ),
	.cout());
defparam \new_state~0 .lut_mask = 16'h8888;
defparam \new_state~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Mux16~0 (
	.dataa(\state[1]~1_combout ),
	.datab(\state[0]~0_combout ),
	.datac(\a_endofpacket~q ),
	.datad(\new_state~0_combout ),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
defparam \Mux16~0 .lut_mask = 16'h06AA;
defparam \Mux16~0 .sum_lutc_input = "datac";

dffeas \state_register[1] (
	.clk(clk),
	.d(\Mux16~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state_register[1]~q ),
	.prn(vcc));
defparam \state_register[1] .is_wysiwyg = "true";
defparam \state_register[1] .power_up = "low";

dffeas \state_d1[1] (
	.clk(clk),
	.d(\state[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state_d1[1]~q ),
	.prn(vcc));
defparam \state_d1[1] .is_wysiwyg = "true";
defparam \state_d1[1] .power_up = "low";

cycloneive_lcell_comb \state[1]~1 (
	.dataa(\state_register[1]~q ),
	.datab(\state_d1[1]~q ),
	.datac(gnd),
	.datad(\in_ready_d1~q ),
	.cin(gnd),
	.combout(\state[1]~1_combout ),
	.cout());
defparam \state[1]~1 .lut_mask = 16'hAACC;
defparam \state[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_valid~0 (
	.dataa(a_valid1),
	.datab(\a_endofpacket~q ),
	.datac(\state[0]~0_combout ),
	.datad(\state[1]~1_combout ),
	.cin(gnd),
	.combout(\out_valid~0_combout ),
	.cout());
defparam \out_valid~0 .lut_mask = 16'hA888;
defparam \out_valid~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \out_valid~1 (
	.dataa(\out_valid~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(a_ready1),
	.cin(gnd),
	.combout(\out_valid~1_combout ),
	.cout());
defparam \out_valid~1 .lut_mask = 16'hAAFF;
defparam \out_valid~1 .sum_lutc_input = "datac";

dffeas \a_data0[0] (
	.clk(clk),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_data0[0]~q ),
	.prn(vcc));
defparam \a_data0[0] .is_wysiwyg = "true";
defparam \a_data0[0] .power_up = "low";

cycloneive_lcell_comb \data0_register[0]~0 (
	.dataa(a_ready1),
	.datab(a_valid1),
	.datac(\state[0]~0_combout ),
	.datad(\state[1]~1_combout ),
	.cin(gnd),
	.combout(\data0_register[0]~0_combout ),
	.cout());
defparam \data0_register[0]~0 .lut_mask = 16'h0008;
defparam \data0_register[0]~0 .sum_lutc_input = "datac";

dffeas \data0_register[0] (
	.clk(clk),
	.d(\a_data0[0]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data0_register[0]~0_combout ),
	.q(\data0_register[0]~q ),
	.prn(vcc));
defparam \data0_register[0] .is_wysiwyg = "true";
defparam \data0_register[0] .power_up = "low";

cycloneive_lcell_comb \b_data[0]~0 (
	.dataa(\data0_register[0]~q ),
	.datab(\a_data0[0]~q ),
	.datac(\state[0]~0_combout ),
	.datad(\state[1]~1_combout ),
	.cin(gnd),
	.combout(\b_data[0]~0_combout ),
	.cout());
defparam \b_data[0]~0 .lut_mask = 16'hAAAC;
defparam \b_data[0]~0 .sum_lutc_input = "datac";

dffeas \a_data0[1] (
	.clk(clk),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_data0[1]~q ),
	.prn(vcc));
defparam \a_data0[1] .is_wysiwyg = "true";
defparam \a_data0[1] .power_up = "low";

dffeas \data0_register[1] (
	.clk(clk),
	.d(\a_data0[1]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data0_register[0]~0_combout ),
	.q(\data0_register[1]~q ),
	.prn(vcc));
defparam \data0_register[1] .is_wysiwyg = "true";
defparam \data0_register[1] .power_up = "low";

cycloneive_lcell_comb \b_data[1]~1 (
	.dataa(\data0_register[1]~q ),
	.datab(\a_data0[1]~q ),
	.datac(\state[0]~0_combout ),
	.datad(\state[1]~1_combout ),
	.cin(gnd),
	.combout(\b_data[1]~1_combout ),
	.cout());
defparam \b_data[1]~1 .lut_mask = 16'hAAAC;
defparam \b_data[1]~1 .sum_lutc_input = "datac";

dffeas \a_data0[2] (
	.clk(clk),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_data0[2]~q ),
	.prn(vcc));
defparam \a_data0[2] .is_wysiwyg = "true";
defparam \a_data0[2] .power_up = "low";

dffeas \data0_register[2] (
	.clk(clk),
	.d(\a_data0[2]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data0_register[0]~0_combout ),
	.q(\data0_register[2]~q ),
	.prn(vcc));
defparam \data0_register[2] .is_wysiwyg = "true";
defparam \data0_register[2] .power_up = "low";

cycloneive_lcell_comb \b_data[2]~2 (
	.dataa(\data0_register[2]~q ),
	.datab(\a_data0[2]~q ),
	.datac(\state[0]~0_combout ),
	.datad(\state[1]~1_combout ),
	.cin(gnd),
	.combout(\b_data[2]~2_combout ),
	.cout());
defparam \b_data[2]~2 .lut_mask = 16'hAAAC;
defparam \b_data[2]~2 .sum_lutc_input = "datac";

dffeas \a_data0[3] (
	.clk(clk),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_data0[3]~q ),
	.prn(vcc));
defparam \a_data0[3] .is_wysiwyg = "true";
defparam \a_data0[3] .power_up = "low";

dffeas \data0_register[3] (
	.clk(clk),
	.d(\a_data0[3]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data0_register[0]~0_combout ),
	.q(\data0_register[3]~q ),
	.prn(vcc));
defparam \data0_register[3] .is_wysiwyg = "true";
defparam \data0_register[3] .power_up = "low";

cycloneive_lcell_comb \b_data[3]~3 (
	.dataa(\data0_register[3]~q ),
	.datab(\a_data0[3]~q ),
	.datac(\state[0]~0_combout ),
	.datad(\state[1]~1_combout ),
	.cin(gnd),
	.combout(\b_data[3]~3_combout ),
	.cout());
defparam \b_data[3]~3 .lut_mask = 16'hAAAC;
defparam \b_data[3]~3 .sum_lutc_input = "datac";

dffeas \a_data0[4] (
	.clk(clk),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_data0[4]~q ),
	.prn(vcc));
defparam \a_data0[4] .is_wysiwyg = "true";
defparam \a_data0[4] .power_up = "low";

dffeas \data0_register[4] (
	.clk(clk),
	.d(\a_data0[4]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data0_register[0]~0_combout ),
	.q(\data0_register[4]~q ),
	.prn(vcc));
defparam \data0_register[4] .is_wysiwyg = "true";
defparam \data0_register[4] .power_up = "low";

cycloneive_lcell_comb \b_data[4]~4 (
	.dataa(\data0_register[4]~q ),
	.datab(\a_data0[4]~q ),
	.datac(\state[0]~0_combout ),
	.datad(\state[1]~1_combout ),
	.cin(gnd),
	.combout(\b_data[4]~4_combout ),
	.cout());
defparam \b_data[4]~4 .lut_mask = 16'hAAAC;
defparam \b_data[4]~4 .sum_lutc_input = "datac";

dffeas \a_data0[5] (
	.clk(clk),
	.d(in_data[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_data0[5]~q ),
	.prn(vcc));
defparam \a_data0[5] .is_wysiwyg = "true";
defparam \a_data0[5] .power_up = "low";

dffeas \data0_register[5] (
	.clk(clk),
	.d(\a_data0[5]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data0_register[0]~0_combout ),
	.q(\data0_register[5]~q ),
	.prn(vcc));
defparam \data0_register[5] .is_wysiwyg = "true";
defparam \data0_register[5] .power_up = "low";

cycloneive_lcell_comb \b_data[5]~5 (
	.dataa(\data0_register[5]~q ),
	.datab(\a_data0[5]~q ),
	.datac(\state[0]~0_combout ),
	.datad(\state[1]~1_combout ),
	.cin(gnd),
	.combout(\b_data[5]~5_combout ),
	.cout());
defparam \b_data[5]~5 .lut_mask = 16'hAAAC;
defparam \b_data[5]~5 .sum_lutc_input = "datac";

dffeas \a_data0[6] (
	.clk(clk),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_data0[6]~q ),
	.prn(vcc));
defparam \a_data0[6] .is_wysiwyg = "true";
defparam \a_data0[6] .power_up = "low";

dffeas \data0_register[6] (
	.clk(clk),
	.d(\a_data0[6]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data0_register[0]~0_combout ),
	.q(\data0_register[6]~q ),
	.prn(vcc));
defparam \data0_register[6] .is_wysiwyg = "true";
defparam \data0_register[6] .power_up = "low";

cycloneive_lcell_comb \b_data[6]~6 (
	.dataa(\data0_register[6]~q ),
	.datab(\a_data0[6]~q ),
	.datac(\state[0]~0_combout ),
	.datad(\state[1]~1_combout ),
	.cin(gnd),
	.combout(\b_data[6]~6_combout ),
	.cout());
defparam \b_data[6]~6 .lut_mask = 16'hAAAC;
defparam \b_data[6]~6 .sum_lutc_input = "datac";

dffeas \a_data0[7] (
	.clk(clk),
	.d(in_data[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_ready1),
	.q(\a_data0[7]~q ),
	.prn(vcc));
defparam \a_data0[7] .is_wysiwyg = "true";
defparam \a_data0[7] .power_up = "low";

dffeas \data0_register[7] (
	.clk(clk),
	.d(\a_data0[7]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data0_register[0]~0_combout ),
	.q(\data0_register[7]~q ),
	.prn(vcc));
defparam \data0_register[7] .is_wysiwyg = "true";
defparam \data0_register[7] .power_up = "low";

cycloneive_lcell_comb \b_data[7]~7 (
	.dataa(\data0_register[7]~q ),
	.datab(\a_data0[7]~q ),
	.datac(\state[0]~0_combout ),
	.datad(\state[1]~1_combout ),
	.cin(gnd),
	.combout(\b_data[7]~7_combout ),
	.cout());
defparam \b_data[7]~7 .lut_mask = 16'hAAAC;
defparam \b_data[7]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \data1_register[0]~0 (
	.dataa(a_ready1),
	.datab(a_valid1),
	.datac(\state[0]~0_combout ),
	.datad(\state[1]~1_combout ),
	.cin(gnd),
	.combout(\data1_register[0]~0_combout ),
	.cout());
defparam \data1_register[0]~0 .lut_mask = 16'h0080;
defparam \data1_register[0]~0 .sum_lutc_input = "datac";

dffeas \data1_register[0] (
	.clk(clk),
	.d(\a_data0[0]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data1_register[0]~0_combout ),
	.q(\data1_register[0]~q ),
	.prn(vcc));
defparam \data1_register[0] .is_wysiwyg = "true";
defparam \data1_register[0] .power_up = "low";

cycloneive_lcell_comb \Mux15~0 (
	.dataa(\data1_register[0]~q ),
	.datab(\state[0]~0_combout ),
	.datac(\a_data0[0]~q ),
	.datad(\state[1]~1_combout ),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
defparam \Mux15~0 .lut_mask = 16'hAAC0;
defparam \Mux15~0 .sum_lutc_input = "datac";

dffeas \data1_register[1] (
	.clk(clk),
	.d(\a_data0[1]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data1_register[0]~0_combout ),
	.q(\data1_register[1]~q ),
	.prn(vcc));
defparam \data1_register[1] .is_wysiwyg = "true";
defparam \data1_register[1] .power_up = "low";

cycloneive_lcell_comb \Mux14~0 (
	.dataa(\data1_register[1]~q ),
	.datab(\state[0]~0_combout ),
	.datac(\a_data0[1]~q ),
	.datad(\state[1]~1_combout ),
	.cin(gnd),
	.combout(\Mux14~0_combout ),
	.cout());
defparam \Mux14~0 .lut_mask = 16'hAAC0;
defparam \Mux14~0 .sum_lutc_input = "datac";

dffeas \data1_register[2] (
	.clk(clk),
	.d(\a_data0[2]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data1_register[0]~0_combout ),
	.q(\data1_register[2]~q ),
	.prn(vcc));
defparam \data1_register[2] .is_wysiwyg = "true";
defparam \data1_register[2] .power_up = "low";

cycloneive_lcell_comb \Mux13~0 (
	.dataa(\data1_register[2]~q ),
	.datab(\state[0]~0_combout ),
	.datac(\a_data0[2]~q ),
	.datad(\state[1]~1_combout ),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
defparam \Mux13~0 .lut_mask = 16'hAAC0;
defparam \Mux13~0 .sum_lutc_input = "datac";

dffeas \data1_register[3] (
	.clk(clk),
	.d(\a_data0[3]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data1_register[0]~0_combout ),
	.q(\data1_register[3]~q ),
	.prn(vcc));
defparam \data1_register[3] .is_wysiwyg = "true";
defparam \data1_register[3] .power_up = "low";

cycloneive_lcell_comb \Mux12~0 (
	.dataa(\data1_register[3]~q ),
	.datab(\state[0]~0_combout ),
	.datac(\a_data0[3]~q ),
	.datad(\state[1]~1_combout ),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
defparam \Mux12~0 .lut_mask = 16'hAAC0;
defparam \Mux12~0 .sum_lutc_input = "datac";

dffeas \data1_register[4] (
	.clk(clk),
	.d(\a_data0[4]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data1_register[0]~0_combout ),
	.q(\data1_register[4]~q ),
	.prn(vcc));
defparam \data1_register[4] .is_wysiwyg = "true";
defparam \data1_register[4] .power_up = "low";

cycloneive_lcell_comb \Mux11~0 (
	.dataa(\data1_register[4]~q ),
	.datab(\state[0]~0_combout ),
	.datac(\a_data0[4]~q ),
	.datad(\state[1]~1_combout ),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
defparam \Mux11~0 .lut_mask = 16'hAAC0;
defparam \Mux11~0 .sum_lutc_input = "datac";

dffeas \data1_register[5] (
	.clk(clk),
	.d(\a_data0[5]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data1_register[0]~0_combout ),
	.q(\data1_register[5]~q ),
	.prn(vcc));
defparam \data1_register[5] .is_wysiwyg = "true";
defparam \data1_register[5] .power_up = "low";

cycloneive_lcell_comb \Mux10~0 (
	.dataa(\data1_register[5]~q ),
	.datab(\state[0]~0_combout ),
	.datac(\a_data0[5]~q ),
	.datad(\state[1]~1_combout ),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
defparam \Mux10~0 .lut_mask = 16'hAAC0;
defparam \Mux10~0 .sum_lutc_input = "datac";

dffeas \data1_register[6] (
	.clk(clk),
	.d(\a_data0[6]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data1_register[0]~0_combout ),
	.q(\data1_register[6]~q ),
	.prn(vcc));
defparam \data1_register[6] .is_wysiwyg = "true";
defparam \data1_register[6] .power_up = "low";

cycloneive_lcell_comb \Mux9~0 (
	.dataa(\data1_register[6]~q ),
	.datab(\state[0]~0_combout ),
	.datac(\a_data0[6]~q ),
	.datad(\state[1]~1_combout ),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
defparam \Mux9~0 .lut_mask = 16'hAAC0;
defparam \Mux9~0 .sum_lutc_input = "datac";

dffeas \data1_register[7] (
	.clk(clk),
	.d(\a_data0[7]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\data1_register[0]~0_combout ),
	.q(\data1_register[7]~q ),
	.prn(vcc));
defparam \data1_register[7] .is_wysiwyg = "true";
defparam \data1_register[7] .power_up = "low";

cycloneive_lcell_comb \Mux8~0 (
	.dataa(\data1_register[7]~q ),
	.datab(\state[0]~0_combout ),
	.datac(\a_data0[7]~q ),
	.datad(\state[1]~1_combout ),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
defparam \Mux8~0 .lut_mask = 16'hAAC0;
defparam \Mux8~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \mem_write2~0 (
	.dataa(a_ready1),
	.datab(a_valid1),
	.datac(\state[1]~1_combout ),
	.datad(\state[0]~0_combout ),
	.cin(gnd),
	.combout(\mem_write2~0_combout ),
	.cout());
defparam \mem_write2~0 .lut_mask = 16'h0080;
defparam \mem_write2~0 .sum_lutc_input = "datac";

dffeas \data2_register[0] (
	.clk(clk),
	.d(\a_data0[0]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_write2~0_combout ),
	.q(\data2_register[0]~q ),
	.prn(vcc));
defparam \data2_register[0] .is_wysiwyg = "true";
defparam \data2_register[0] .power_up = "low";

cycloneive_lcell_comb \Mux7~0 (
	.dataa(\state[1]~1_combout ),
	.datab(\data2_register[0]~q ),
	.datac(\a_data0[0]~q ),
	.datad(\state[0]~0_combout ),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
defparam \Mux7~0 .lut_mask = 16'h88A0;
defparam \Mux7~0 .sum_lutc_input = "datac";

dffeas \data2_register[1] (
	.clk(clk),
	.d(\a_data0[1]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_write2~0_combout ),
	.q(\data2_register[1]~q ),
	.prn(vcc));
defparam \data2_register[1] .is_wysiwyg = "true";
defparam \data2_register[1] .power_up = "low";

cycloneive_lcell_comb \Mux6~0 (
	.dataa(\state[1]~1_combout ),
	.datab(\data2_register[1]~q ),
	.datac(\a_data0[1]~q ),
	.datad(\state[0]~0_combout ),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
defparam \Mux6~0 .lut_mask = 16'h88A0;
defparam \Mux6~0 .sum_lutc_input = "datac";

dffeas \data2_register[2] (
	.clk(clk),
	.d(\a_data0[2]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_write2~0_combout ),
	.q(\data2_register[2]~q ),
	.prn(vcc));
defparam \data2_register[2] .is_wysiwyg = "true";
defparam \data2_register[2] .power_up = "low";

cycloneive_lcell_comb \Mux5~0 (
	.dataa(\state[1]~1_combout ),
	.datab(\data2_register[2]~q ),
	.datac(\a_data0[2]~q ),
	.datad(\state[0]~0_combout ),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
defparam \Mux5~0 .lut_mask = 16'h88A0;
defparam \Mux5~0 .sum_lutc_input = "datac";

dffeas \data2_register[3] (
	.clk(clk),
	.d(\a_data0[3]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_write2~0_combout ),
	.q(\data2_register[3]~q ),
	.prn(vcc));
defparam \data2_register[3] .is_wysiwyg = "true";
defparam \data2_register[3] .power_up = "low";

cycloneive_lcell_comb \Mux4~0 (
	.dataa(\state[1]~1_combout ),
	.datab(\data2_register[3]~q ),
	.datac(\a_data0[3]~q ),
	.datad(\state[0]~0_combout ),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
defparam \Mux4~0 .lut_mask = 16'h88A0;
defparam \Mux4~0 .sum_lutc_input = "datac";

dffeas \data2_register[4] (
	.clk(clk),
	.d(\a_data0[4]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_write2~0_combout ),
	.q(\data2_register[4]~q ),
	.prn(vcc));
defparam \data2_register[4] .is_wysiwyg = "true";
defparam \data2_register[4] .power_up = "low";

cycloneive_lcell_comb \Mux3~0 (
	.dataa(\state[1]~1_combout ),
	.datab(\data2_register[4]~q ),
	.datac(\a_data0[4]~q ),
	.datad(\state[0]~0_combout ),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
defparam \Mux3~0 .lut_mask = 16'h88A0;
defparam \Mux3~0 .sum_lutc_input = "datac";

dffeas \data2_register[5] (
	.clk(clk),
	.d(\a_data0[5]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_write2~0_combout ),
	.q(\data2_register[5]~q ),
	.prn(vcc));
defparam \data2_register[5] .is_wysiwyg = "true";
defparam \data2_register[5] .power_up = "low";

cycloneive_lcell_comb \Mux2~0 (
	.dataa(\state[1]~1_combout ),
	.datab(\data2_register[5]~q ),
	.datac(\a_data0[5]~q ),
	.datad(\state[0]~0_combout ),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
defparam \Mux2~0 .lut_mask = 16'h88A0;
defparam \Mux2~0 .sum_lutc_input = "datac";

dffeas \data2_register[6] (
	.clk(clk),
	.d(\a_data0[6]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_write2~0_combout ),
	.q(\data2_register[6]~q ),
	.prn(vcc));
defparam \data2_register[6] .is_wysiwyg = "true";
defparam \data2_register[6] .power_up = "low";

cycloneive_lcell_comb \Mux1~0 (
	.dataa(\state[1]~1_combout ),
	.datab(\data2_register[6]~q ),
	.datac(\a_data0[6]~q ),
	.datad(\state[0]~0_combout ),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
defparam \Mux1~0 .lut_mask = 16'h88A0;
defparam \Mux1~0 .sum_lutc_input = "datac";

dffeas \data2_register[7] (
	.clk(clk),
	.d(\a_data0[7]~q ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_write2~0_combout ),
	.q(\data2_register[7]~q ),
	.prn(vcc));
defparam \data2_register[7] .is_wysiwyg = "true";
defparam \data2_register[7] .power_up = "low";

cycloneive_lcell_comb \Mux0~0 (
	.dataa(\state[1]~1_combout ),
	.datab(\data2_register[7]~q ),
	.datac(\a_data0[7]~q ),
	.datad(\state[0]~0_combout ),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'h88A0;
defparam \Mux0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_data[24]~8 (
	.dataa(\state[0]~0_combout ),
	.datab(\state[1]~1_combout ),
	.datac(\a_data0[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\b_data[24]~8_combout ),
	.cout());
defparam \b_data[24]~8 .lut_mask = 16'h8080;
defparam \b_data[24]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_data[25]~9 (
	.dataa(\state[0]~0_combout ),
	.datab(\state[1]~1_combout ),
	.datac(\a_data0[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\b_data[25]~9_combout ),
	.cout());
defparam \b_data[25]~9 .lut_mask = 16'h8080;
defparam \b_data[25]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_data[26]~10 (
	.dataa(\state[0]~0_combout ),
	.datab(\state[1]~1_combout ),
	.datac(\a_data0[2]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\b_data[26]~10_combout ),
	.cout());
defparam \b_data[26]~10 .lut_mask = 16'h8080;
defparam \b_data[26]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_data[27]~11 (
	.dataa(\state[0]~0_combout ),
	.datab(\state[1]~1_combout ),
	.datac(\a_data0[3]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\b_data[27]~11_combout ),
	.cout());
defparam \b_data[27]~11 .lut_mask = 16'h8080;
defparam \b_data[27]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_data[28]~12 (
	.dataa(\state[0]~0_combout ),
	.datab(\state[1]~1_combout ),
	.datac(\a_data0[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\b_data[28]~12_combout ),
	.cout());
defparam \b_data[28]~12 .lut_mask = 16'h8080;
defparam \b_data[28]~12 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_data[29]~13 (
	.dataa(\state[0]~0_combout ),
	.datab(\state[1]~1_combout ),
	.datac(\a_data0[5]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\b_data[29]~13_combout ),
	.cout());
defparam \b_data[29]~13 .lut_mask = 16'h8080;
defparam \b_data[29]~13 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_data[30]~14 (
	.dataa(\state[0]~0_combout ),
	.datab(\state[1]~1_combout ),
	.datac(\a_data0[6]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\b_data[30]~14_combout ),
	.cout());
defparam \b_data[30]~14 .lut_mask = 16'h8080;
defparam \b_data[30]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \b_data[31]~15 (
	.dataa(\state[0]~0_combout ),
	.datab(\state[1]~1_combout ),
	.datac(\a_data0[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\b_data[31]~15_combout ),
	.cout());
defparam \b_data[31]~15 .lut_mask = 16'h8080;
defparam \b_data[31]~15 .sum_lutc_input = "datac";

endmodule

module flashLoader_intel_generic_serial_flash_interface_csr (
	avl_rddata_local_0,
	avl_rddata_local_1,
	avl_rddata_local_2,
	avl_rddata_local_3,
	avl_rddata_local_4,
	avl_rddata_local_5,
	avl_rddata_local_6,
	avl_rddata_local_7,
	avl_rddata_local_8,
	avl_rddata_local_9,
	avl_rddata_local_10,
	avl_rddata_local_11,
	avl_rddata_local_12,
	avl_rddata_local_13,
	avl_rddata_local_14,
	avl_rddata_local_15,
	avl_rddata_local_16,
	avl_rddata_local_17,
	avl_rddata_local_18,
	avl_rddata_local_19,
	avl_rddata_local_20,
	avl_rddata_local_21,
	avl_rddata_local_22,
	avl_rddata_local_23,
	avl_rddata_local_24,
	avl_rddata_local_25,
	avl_rddata_local_26,
	avl_rddata_local_27,
	avl_rddata_local_28,
	avl_rddata_local_29,
	avl_rddata_local_30,
	avl_rddata_local_31,
	stateST_IDLE,
	hold_waitrequest,
	csr_waitrequest1,
	avl_rddatavalid_local1,
	csr_wr_inst_data_0,
	csr_rd_inst_data_0,
	csr_op_protocol_data_0,
	csr_flash_cmd_wr_data_0_data_0,
	csr_flash_cmd_addr_data_0,
	csr_flash_cmd_wr_data_1_data_0,
	csr_delay_setting_data_0,
	csr_clk_baud_rate_data_0,
	csr_control_data_0,
	csr_rd_capturing_data_0,
	reset,
	csr_wr_inst_data_1,
	csr_rd_inst_data_1,
	csr_op_protocol_data_1,
	csr_flash_cmd_wr_data_0_data_1,
	csr_flash_cmd_addr_data_1,
	csr_flash_cmd_wr_data_1_data_1,
	csr_delay_setting_data_1,
	csr_clk_baud_rate_data_1,
	csr_rd_capturing_data_1,
	csr_wr_inst_data_2,
	csr_rd_inst_data_2,
	csr_flash_cmd_wr_data_0_data_2,
	csr_flash_cmd_addr_data_2,
	csr_flash_cmd_wr_data_1_data_2,
	csr_delay_setting_data_2,
	csr_clk_baud_rate_data_2,
	csr_rd_capturing_data_2,
	csr_wr_inst_data_3,
	csr_rd_inst_data_3,
	csr_flash_cmd_wr_data_0_data_3,
	csr_flash_cmd_addr_data_3,
	csr_flash_cmd_wr_data_1_data_3,
	csr_delay_setting_data_3,
	csr_clk_baud_rate_data_3,
	csr_rd_capturing_data_3,
	csr_wr_inst_data_4,
	csr_delay_setting_data_4,
	csr_flash_cmd_addr_data_4,
	csr_op_protocol_data_4,
	csr_clk_baud_rate_data_4,
	csr_control_data_4,
	csr_rd_inst_data_4,
	csr_flash_cmd_wr_data_1_data_4,
	csr_flash_cmd_wr_data_0_data_4,
	csr_delay_setting_data_5,
	csr_wr_inst_data_5,
	csr_rd_inst_data_5,
	csr_op_protocol_data_5,
	csr_control_data_5,
	csr_flash_cmd_wr_data_1_data_5,
	csr_flash_cmd_wr_data_0_data_5,
	csr_flash_cmd_addr_data_5,
	csr_wr_inst_data_6,
	csr_rd_inst_data_6,
	csr_delay_setting_data_6,
	csr_control_data_6,
	csr_flash_cmd_wr_data_1_data_6,
	csr_flash_cmd_wr_data_0_data_6,
	csr_flash_cmd_addr_data_6,
	csr_delay_setting_data_7,
	csr_wr_inst_data_7,
	csr_rd_inst_data_7,
	csr_control_data_7,
	csr_flash_cmd_wr_data_1_data_7,
	csr_flash_cmd_wr_data_0_data_7,
	csr_flash_cmd_addr_data_7,
	csr_rd_inst_data_8,
	csr_op_protocol_data_8,
	csr_flash_cmd_addr_data_8,
	csr_control_data_8,
	csr_flash_cmd_wr_data_0_data_8,
	csr_wr_inst_data_8,
	csr_flash_cmd_wr_data_1_data_8,
	csr_flash_cmd_addr_data_9,
	csr_rd_inst_data_9,
	csr_op_protocol_data_9,
	csr_flash_cmd_wr_data_0_data_9,
	csr_wr_inst_data_9,
	csr_flash_cmd_wr_data_1_data_9,
	csr_rd_inst_data_10,
	csr_flash_cmd_addr_data_10,
	csr_flash_cmd_wr_data_0_data_10,
	csr_wr_inst_data_10,
	csr_flash_cmd_wr_data_1_data_10,
	csr_flash_cmd_addr_data_11,
	csr_rd_inst_data_11,
	csr_flash_cmd_wr_data_0_data_11,
	csr_wr_inst_data_11,
	csr_flash_cmd_wr_data_1_data_11,
	csr_rd_inst_data_12,
	csr_op_protocol_data_12,
	csr_flash_cmd_addr_data_12,
	csr_flash_cmd_wr_data_0_data_12,
	csr_wr_inst_data_12,
	csr_flash_cmd_wr_data_1_data_12,
	csr_flash_cmd_addr_data_13,
	csr_op_protocol_data_13,
	csr_flash_cmd_wr_data_0_data_13,
	csr_wr_inst_data_13,
	csr_flash_cmd_wr_data_1_data_13,
	csr_flash_cmd_addr_data_14,
	csr_flash_cmd_wr_data_0_data_14,
	csr_wr_inst_data_14,
	csr_flash_cmd_wr_data_1_data_14,
	csr_flash_cmd_addr_data_15,
	csr_flash_cmd_wr_data_0_data_15,
	csr_wr_inst_data_15,
	csr_flash_cmd_wr_data_1_data_15,
	csr_op_protocol_data_16,
	csr_flash_cmd_addr_data_16,
	csr_flash_cmd_wr_data_0_data_16,
	csr_flash_cmd_wr_data_1_data_16,
	csr_flash_cmd_addr_data_17,
	csr_op_protocol_data_17,
	csr_flash_cmd_wr_data_0_data_17,
	csr_flash_cmd_wr_data_1_data_17,
	csr_flash_cmd_addr_data_18,
	csr_flash_cmd_wr_data_0_data_18,
	csr_flash_cmd_wr_data_1_data_18,
	csr_flash_cmd_addr_data_19,
	csr_flash_cmd_wr_data_0_data_19,
	csr_flash_cmd_wr_data_1_data_19,
	csr_flash_cmd_addr_data_20,
	csr_flash_cmd_wr_data_0_data_20,
	csr_flash_cmd_wr_data_1_data_20,
	csr_flash_cmd_addr_data_21,
	csr_flash_cmd_wr_data_0_data_21,
	csr_flash_cmd_wr_data_1_data_21,
	csr_flash_cmd_addr_data_22,
	csr_flash_cmd_wr_data_0_data_22,
	csr_flash_cmd_wr_data_1_data_22,
	csr_flash_cmd_addr_data_23,
	csr_flash_cmd_wr_data_0_data_23,
	csr_flash_cmd_wr_data_1_data_23,
	csr_flash_cmd_addr_data_24,
	csr_flash_cmd_wr_data_0_data_24,
	csr_flash_cmd_wr_data_1_data_24,
	csr_flash_cmd_addr_data_25,
	csr_flash_cmd_wr_data_0_data_25,
	csr_flash_cmd_wr_data_1_data_25,
	csr_flash_cmd_addr_data_26,
	csr_flash_cmd_wr_data_0_data_26,
	csr_flash_cmd_wr_data_1_data_26,
	csr_flash_cmd_addr_data_27,
	csr_flash_cmd_wr_data_0_data_27,
	csr_flash_cmd_wr_data_1_data_27,
	csr_flash_cmd_addr_data_28,
	csr_flash_cmd_wr_data_0_data_28,
	csr_flash_cmd_wr_data_1_data_28,
	csr_flash_cmd_addr_data_29,
	csr_flash_cmd_wr_data_0_data_29,
	csr_flash_cmd_wr_data_1_data_29,
	csr_flash_cmd_addr_data_30,
	csr_flash_cmd_wr_data_0_data_30,
	csr_flash_cmd_wr_data_1_data_30,
	csr_flash_cmd_addr_data_31,
	csr_flash_cmd_wr_data_0_data_31,
	csr_flash_cmd_wr_data_1_data_31,
	stateST_SEND_DUMMY_RSP,
	out_valid,
	out_endofpacket,
	in_cmd_channel_reg_1,
	stateST_WAIT_RSP,
	sink_ready,
	out_rsp_data_0,
	out_rsp_data_1,
	out_rsp_data_2,
	out_rsp_data_3,
	out_rsp_data_4,
	out_rsp_data_5,
	out_rsp_data_6,
	out_rsp_data_7,
	out_rsp_data_8,
	out_rsp_data_9,
	out_rsp_data_10,
	out_rsp_data_11,
	out_rsp_data_12,
	out_rsp_data_13,
	out_rsp_data_14,
	out_rsp_data_15,
	out_rsp_data_16,
	out_rsp_data_17,
	out_rsp_data_18,
	out_rsp_data_19,
	out_rsp_data_20,
	out_rsp_data_21,
	out_rsp_data_22,
	out_rsp_data_23,
	out_rsp_data_24,
	out_rsp_data_25,
	out_rsp_data_26,
	out_rsp_data_27,
	out_rsp_data_28,
	out_rsp_data_29,
	out_rsp_data_30,
	out_rsp_data_31,
	saved_grant_1,
	stateST_SEND_HEADER,
	stateST_SEND_DATA_1,
	stateST_SEND_DATA_0,
	has_data_in1,
	more_than_4bytes_data1,
	src_payload_0,
	Selector18,
	sink1_ready,
	Selector34,
	has_data_out1,
	numb_data_0,
	numb_data_1,
	numb_data_3,
	numb_data_2,
	has_addr1,
	numb_dummy_0,
	numb_dummy_4,
	numb_dummy_3,
	numb_dummy_2,
	numb_dummy_1,
	is_4bytes_addr1,
	opcode_0,
	opcode_4,
	opcode_2,
	opcode_1,
	opcode_3,
	opcode_5,
	opcode_6,
	opcode_7,
	has_dummy1,
	avl_csr_address_1,
	avl_csr_address_0,
	avl_csr_address_2,
	avl_csr_address_3,
	avl_csr_read,
	avl_csr_address_4,
	avl_csr_address_5,
	clk,
	avl_csr_write,
	csr_wrdata)/* synthesis synthesis_greybox=0 */;
output 	avl_rddata_local_0;
output 	avl_rddata_local_1;
output 	avl_rddata_local_2;
output 	avl_rddata_local_3;
output 	avl_rddata_local_4;
output 	avl_rddata_local_5;
output 	avl_rddata_local_6;
output 	avl_rddata_local_7;
output 	avl_rddata_local_8;
output 	avl_rddata_local_9;
output 	avl_rddata_local_10;
output 	avl_rddata_local_11;
output 	avl_rddata_local_12;
output 	avl_rddata_local_13;
output 	avl_rddata_local_14;
output 	avl_rddata_local_15;
output 	avl_rddata_local_16;
output 	avl_rddata_local_17;
output 	avl_rddata_local_18;
output 	avl_rddata_local_19;
output 	avl_rddata_local_20;
output 	avl_rddata_local_21;
output 	avl_rddata_local_22;
output 	avl_rddata_local_23;
output 	avl_rddata_local_24;
output 	avl_rddata_local_25;
output 	avl_rddata_local_26;
output 	avl_rddata_local_27;
output 	avl_rddata_local_28;
output 	avl_rddata_local_29;
output 	avl_rddata_local_30;
output 	avl_rddata_local_31;
output 	stateST_IDLE;
input 	hold_waitrequest;
output 	csr_waitrequest1;
output 	avl_rddatavalid_local1;
output 	csr_wr_inst_data_0;
output 	csr_rd_inst_data_0;
output 	csr_op_protocol_data_0;
output 	csr_flash_cmd_wr_data_0_data_0;
output 	csr_flash_cmd_addr_data_0;
output 	csr_flash_cmd_wr_data_1_data_0;
output 	csr_delay_setting_data_0;
output 	csr_clk_baud_rate_data_0;
output 	csr_control_data_0;
output 	csr_rd_capturing_data_0;
input 	reset;
output 	csr_wr_inst_data_1;
output 	csr_rd_inst_data_1;
output 	csr_op_protocol_data_1;
output 	csr_flash_cmd_wr_data_0_data_1;
output 	csr_flash_cmd_addr_data_1;
output 	csr_flash_cmd_wr_data_1_data_1;
output 	csr_delay_setting_data_1;
output 	csr_clk_baud_rate_data_1;
output 	csr_rd_capturing_data_1;
output 	csr_wr_inst_data_2;
output 	csr_rd_inst_data_2;
output 	csr_flash_cmd_wr_data_0_data_2;
output 	csr_flash_cmd_addr_data_2;
output 	csr_flash_cmd_wr_data_1_data_2;
output 	csr_delay_setting_data_2;
output 	csr_clk_baud_rate_data_2;
output 	csr_rd_capturing_data_2;
output 	csr_wr_inst_data_3;
output 	csr_rd_inst_data_3;
output 	csr_flash_cmd_wr_data_0_data_3;
output 	csr_flash_cmd_addr_data_3;
output 	csr_flash_cmd_wr_data_1_data_3;
output 	csr_delay_setting_data_3;
output 	csr_clk_baud_rate_data_3;
output 	csr_rd_capturing_data_3;
output 	csr_wr_inst_data_4;
output 	csr_delay_setting_data_4;
output 	csr_flash_cmd_addr_data_4;
output 	csr_op_protocol_data_4;
output 	csr_clk_baud_rate_data_4;
output 	csr_control_data_4;
output 	csr_rd_inst_data_4;
output 	csr_flash_cmd_wr_data_1_data_4;
output 	csr_flash_cmd_wr_data_0_data_4;
output 	csr_delay_setting_data_5;
output 	csr_wr_inst_data_5;
output 	csr_rd_inst_data_5;
output 	csr_op_protocol_data_5;
output 	csr_control_data_5;
output 	csr_flash_cmd_wr_data_1_data_5;
output 	csr_flash_cmd_wr_data_0_data_5;
output 	csr_flash_cmd_addr_data_5;
output 	csr_wr_inst_data_6;
output 	csr_rd_inst_data_6;
output 	csr_delay_setting_data_6;
output 	csr_control_data_6;
output 	csr_flash_cmd_wr_data_1_data_6;
output 	csr_flash_cmd_wr_data_0_data_6;
output 	csr_flash_cmd_addr_data_6;
output 	csr_delay_setting_data_7;
output 	csr_wr_inst_data_7;
output 	csr_rd_inst_data_7;
output 	csr_control_data_7;
output 	csr_flash_cmd_wr_data_1_data_7;
output 	csr_flash_cmd_wr_data_0_data_7;
output 	csr_flash_cmd_addr_data_7;
output 	csr_rd_inst_data_8;
output 	csr_op_protocol_data_8;
output 	csr_flash_cmd_addr_data_8;
output 	csr_control_data_8;
output 	csr_flash_cmd_wr_data_0_data_8;
output 	csr_wr_inst_data_8;
output 	csr_flash_cmd_wr_data_1_data_8;
output 	csr_flash_cmd_addr_data_9;
output 	csr_rd_inst_data_9;
output 	csr_op_protocol_data_9;
output 	csr_flash_cmd_wr_data_0_data_9;
output 	csr_wr_inst_data_9;
output 	csr_flash_cmd_wr_data_1_data_9;
output 	csr_rd_inst_data_10;
output 	csr_flash_cmd_addr_data_10;
output 	csr_flash_cmd_wr_data_0_data_10;
output 	csr_wr_inst_data_10;
output 	csr_flash_cmd_wr_data_1_data_10;
output 	csr_flash_cmd_addr_data_11;
output 	csr_rd_inst_data_11;
output 	csr_flash_cmd_wr_data_0_data_11;
output 	csr_wr_inst_data_11;
output 	csr_flash_cmd_wr_data_1_data_11;
output 	csr_rd_inst_data_12;
output 	csr_op_protocol_data_12;
output 	csr_flash_cmd_addr_data_12;
output 	csr_flash_cmd_wr_data_0_data_12;
output 	csr_wr_inst_data_12;
output 	csr_flash_cmd_wr_data_1_data_12;
output 	csr_flash_cmd_addr_data_13;
output 	csr_op_protocol_data_13;
output 	csr_flash_cmd_wr_data_0_data_13;
output 	csr_wr_inst_data_13;
output 	csr_flash_cmd_wr_data_1_data_13;
output 	csr_flash_cmd_addr_data_14;
output 	csr_flash_cmd_wr_data_0_data_14;
output 	csr_wr_inst_data_14;
output 	csr_flash_cmd_wr_data_1_data_14;
output 	csr_flash_cmd_addr_data_15;
output 	csr_flash_cmd_wr_data_0_data_15;
output 	csr_wr_inst_data_15;
output 	csr_flash_cmd_wr_data_1_data_15;
output 	csr_op_protocol_data_16;
output 	csr_flash_cmd_addr_data_16;
output 	csr_flash_cmd_wr_data_0_data_16;
output 	csr_flash_cmd_wr_data_1_data_16;
output 	csr_flash_cmd_addr_data_17;
output 	csr_op_protocol_data_17;
output 	csr_flash_cmd_wr_data_0_data_17;
output 	csr_flash_cmd_wr_data_1_data_17;
output 	csr_flash_cmd_addr_data_18;
output 	csr_flash_cmd_wr_data_0_data_18;
output 	csr_flash_cmd_wr_data_1_data_18;
output 	csr_flash_cmd_addr_data_19;
output 	csr_flash_cmd_wr_data_0_data_19;
output 	csr_flash_cmd_wr_data_1_data_19;
output 	csr_flash_cmd_addr_data_20;
output 	csr_flash_cmd_wr_data_0_data_20;
output 	csr_flash_cmd_wr_data_1_data_20;
output 	csr_flash_cmd_addr_data_21;
output 	csr_flash_cmd_wr_data_0_data_21;
output 	csr_flash_cmd_wr_data_1_data_21;
output 	csr_flash_cmd_addr_data_22;
output 	csr_flash_cmd_wr_data_0_data_22;
output 	csr_flash_cmd_wr_data_1_data_22;
output 	csr_flash_cmd_addr_data_23;
output 	csr_flash_cmd_wr_data_0_data_23;
output 	csr_flash_cmd_wr_data_1_data_23;
output 	csr_flash_cmd_addr_data_24;
output 	csr_flash_cmd_wr_data_0_data_24;
output 	csr_flash_cmd_wr_data_1_data_24;
output 	csr_flash_cmd_addr_data_25;
output 	csr_flash_cmd_wr_data_0_data_25;
output 	csr_flash_cmd_wr_data_1_data_25;
output 	csr_flash_cmd_addr_data_26;
output 	csr_flash_cmd_wr_data_0_data_26;
output 	csr_flash_cmd_wr_data_1_data_26;
output 	csr_flash_cmd_addr_data_27;
output 	csr_flash_cmd_wr_data_0_data_27;
output 	csr_flash_cmd_wr_data_1_data_27;
output 	csr_flash_cmd_addr_data_28;
output 	csr_flash_cmd_wr_data_0_data_28;
output 	csr_flash_cmd_wr_data_1_data_28;
output 	csr_flash_cmd_addr_data_29;
output 	csr_flash_cmd_wr_data_0_data_29;
output 	csr_flash_cmd_wr_data_1_data_29;
output 	csr_flash_cmd_addr_data_30;
output 	csr_flash_cmd_wr_data_0_data_30;
output 	csr_flash_cmd_wr_data_1_data_30;
output 	csr_flash_cmd_addr_data_31;
output 	csr_flash_cmd_wr_data_0_data_31;
output 	csr_flash_cmd_wr_data_1_data_31;
input 	stateST_SEND_DUMMY_RSP;
input 	out_valid;
input 	out_endofpacket;
input 	in_cmd_channel_reg_1;
output 	stateST_WAIT_RSP;
input 	sink_ready;
input 	out_rsp_data_0;
input 	out_rsp_data_1;
input 	out_rsp_data_2;
input 	out_rsp_data_3;
input 	out_rsp_data_4;
input 	out_rsp_data_5;
input 	out_rsp_data_6;
input 	out_rsp_data_7;
input 	out_rsp_data_8;
input 	out_rsp_data_9;
input 	out_rsp_data_10;
input 	out_rsp_data_11;
input 	out_rsp_data_12;
input 	out_rsp_data_13;
input 	out_rsp_data_14;
input 	out_rsp_data_15;
input 	out_rsp_data_16;
input 	out_rsp_data_17;
input 	out_rsp_data_18;
input 	out_rsp_data_19;
input 	out_rsp_data_20;
input 	out_rsp_data_21;
input 	out_rsp_data_22;
input 	out_rsp_data_23;
input 	out_rsp_data_24;
input 	out_rsp_data_25;
input 	out_rsp_data_26;
input 	out_rsp_data_27;
input 	out_rsp_data_28;
input 	out_rsp_data_29;
input 	out_rsp_data_30;
input 	out_rsp_data_31;
input 	saved_grant_1;
output 	stateST_SEND_HEADER;
output 	stateST_SEND_DATA_1;
output 	stateST_SEND_DATA_0;
output 	has_data_in1;
output 	more_than_4bytes_data1;
input 	src_payload_0;
input 	Selector18;
input 	sink1_ready;
output 	Selector34;
output 	has_data_out1;
output 	numb_data_0;
output 	numb_data_1;
output 	numb_data_3;
output 	numb_data_2;
output 	has_addr1;
output 	numb_dummy_0;
output 	numb_dummy_4;
output 	numb_dummy_3;
output 	numb_dummy_2;
output 	numb_dummy_1;
output 	is_4bytes_addr1;
output 	opcode_0;
output 	opcode_4;
output 	opcode_2;
output 	opcode_1;
output 	opcode_3;
output 	opcode_5;
output 	opcode_6;
output 	opcode_7;
output 	has_dummy1;
input 	avl_csr_address_1;
input 	avl_csr_address_0;
input 	avl_csr_address_2;
input 	avl_csr_address_3;
input 	avl_csr_read;
input 	avl_csr_address_4;
input 	avl_csr_address_5;
input 	clk;
input 	avl_csr_write;
input 	[31:0] csr_wrdata;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \rdata_comb[0]~2_combout ;
wire \csr_flash_cmd_setting_data[0]~0_combout ;
wire \wr_csr_control~0_combout ;
wire \wr_csr_op_protocol~0_combout ;
wire \wr_csr_flash_cmd_setting~combout ;
wire \csr_flash_cmd_setting_data[0]~q ;
wire \rdata_comb[0]~3_combout ;
wire \avl_rddata_local[3]~2_combout ;
wire \avl_rddata_local[3]~3_combout ;
wire \read_data_cnt~1_combout ;
wire \read_data_cnt[0]~2_combout ;
wire \read_data_cnt[0]~q ;
wire \read_data_cnt~3_combout ;
wire \read_data_cnt[1]~q ;
wire \csr_flash_cmd_rd_data_0_data[0]~0_combout ;
wire \csr_flash_cmd_rd_data_0_data[0]~q ;
wire \avl_rddata_local[3]~4_combout ;
wire \rdata_comb[0]~4_combout ;
wire \rdata_comb[0]~5_combout ;
wire \rdata_comb[0]~6_combout ;
wire \rdata_comb[0]~7_combout ;
wire \rdata_comb[0]~8_combout ;
wire \csr_flash_cmd_rd_data_1_data[0]~0_combout ;
wire \csr_flash_cmd_rd_data_1_data[0]~q ;
wire \rdata_comb[0]~9_combout ;
wire \rdata_comb[4]~10_combout ;
wire \avl_rddata_local[3]~5_combout ;
wire \rdata_comb[0]~11_combout ;
wire \rdata_comb[1]~12_combout ;
wire \csr_flash_cmd_setting_data[1]~q ;
wire \rdata_comb[1]~13_combout ;
wire \csr_flash_cmd_rd_data_0_data[1]~q ;
wire \rdata_comb[1]~14_combout ;
wire \rdata_comb[1]~15_combout ;
wire \wr_csr_control~1_combout ;
wire \wr_csr_control~combout ;
wire \csr_control_data[1]~q ;
wire \rdata_comb[1]~16_combout ;
wire \rdata_comb[1]~17_combout ;
wire \rdata_comb[1]~18_combout ;
wire \csr_flash_cmd_rd_data_1_data[1]~q ;
wire \rdata_comb[1]~19_combout ;
wire \rdata_comb[1]~20_combout ;
wire \wr_csr_op_protocol~combout ;
wire \csr_op_protocol_data[2]~q ;
wire \rdata_comb[2]~21_combout ;
wire \csr_flash_cmd_setting_data[2]~1_combout ;
wire \csr_flash_cmd_setting_data[2]~q ;
wire \rdata_comb[2]~22_combout ;
wire \csr_flash_cmd_rd_data_0_data[2]~q ;
wire \rdata_comb[2]~23_combout ;
wire \rdata_comb[2]~24_combout ;
wire \csr_control_data[2]~q ;
wire \rdata_comb[2]~25_combout ;
wire \rdata_comb[2]~26_combout ;
wire \rdata_comb[2]~27_combout ;
wire \csr_flash_cmd_rd_data_1_data[2]~q ;
wire \rdata_comb[2]~28_combout ;
wire \rdata_comb[2]~29_combout ;
wire \csr_op_protocol_data[3]~q ;
wire \rdata_comb[3]~30_combout ;
wire \csr_flash_cmd_setting_data[3]~q ;
wire \rdata_comb[3]~31_combout ;
wire \csr_flash_cmd_rd_data_0_data[3]~q ;
wire \rdata_comb[3]~32_combout ;
wire \rdata_comb[3]~33_combout ;
wire \csr_control_data[3]~q ;
wire \rdata_comb[3]~34_combout ;
wire \rdata_comb[3]~35_combout ;
wire \rdata_comb[3]~36_combout ;
wire \csr_flash_cmd_rd_data_1_data[3]~q ;
wire \rdata_comb[3]~37_combout ;
wire \rdata_comb[3]~38_combout ;
wire \Selector27~0_combout ;
wire \csr_flash_cmd_setting_data[4]~q ;
wire \Selector27~1_combout ;
wire \csr_flash_cmd_rd_data_1_data[4]~q ;
wire \csr_flash_cmd_rd_data_0_data[4]~q ;
wire \Selector27~2_combout ;
wire \Selector27~3_combout ;
wire \Selector27~4_combout ;
wire \Selector27~5_combout ;
wire \Selector27~6_combout ;
wire \Selector27~7_combout ;
wire \Selector27~8_combout ;
wire \rdata_comb[4]~235_combout ;
wire \wr_csr_flash_cmd_addr~0_combout ;
wire \csr_flash_cmd_rd_data_1_data[5]~q ;
wire \rdata_comb[5]~39_combout ;
wire \avl_rddata_local[7]~6_combout ;
wire \rdata_comb[5]~40_combout ;
wire \csr_flash_cmd_setting_data[5]~q ;
wire \rdata_comb[5]~41_combout ;
wire \avl_rddata_local[7]~7_combout ;
wire \rdata_comb[5]~42_combout ;
wire \csr_flash_cmd_rd_data_0_data[5]~q ;
wire \rdata_comb[5]~43_combout ;
wire \rdata_comb[5]~44_combout ;
wire \rdata_comb[5]~45_combout ;
wire \rdata_comb[5]~46_combout ;
wire \rdata_comb[5]~47_combout ;
wire \rdata_comb[5]~48_combout ;
wire \csr_flash_cmd_rd_data_1_data[6]~q ;
wire \rdata_comb[6]~49_combout ;
wire \csr_op_protocol_data[6]~q ;
wire \rdata_comb[6]~50_combout ;
wire \csr_flash_cmd_setting_data[6]~q ;
wire \rdata_comb[6]~51_combout ;
wire \rdata_comb[6]~52_combout ;
wire \csr_flash_cmd_rd_data_0_data[6]~q ;
wire \rdata_comb[6]~53_combout ;
wire \rdata_comb[6]~54_combout ;
wire \rdata_comb[6]~55_combout ;
wire \rdata_comb[6]~56_combout ;
wire \rdata_comb[6]~57_combout ;
wire \csr_flash_cmd_rd_data_1_data[7]~q ;
wire \rdata_comb[7]~58_combout ;
wire \csr_op_protocol_data[7]~q ;
wire \rdata_comb[7]~59_combout ;
wire \csr_flash_cmd_setting_data[7]~q ;
wire \rdata_comb[7]~60_combout ;
wire \rdata_comb[7]~61_combout ;
wire \csr_flash_cmd_rd_data_0_data[7]~q ;
wire \rdata_comb[7]~62_combout ;
wire \rdata_comb[7]~63_combout ;
wire \rdata_comb[7]~64_combout ;
wire \rdata_comb[7]~65_combout ;
wire \rdata_comb[7]~66_combout ;
wire \csr_flash_cmd_rd_data_0_data[8]~q ;
wire \rdata_comb[8]~67_combout ;
wire \csr_flash_cmd_rd_data_1_data[8]~q ;
wire \rdata_comb[8]~68_combout ;
wire \avl_rddata_local[13]~8_combout ;
wire \avl_rddata_local[13]~9_combout ;
wire \rdata_comb[8]~69_combout ;
wire \csr_flash_cmd_setting_data[8]~q ;
wire \rdata_comb[8]~70_combout ;
wire \rdata_comb[8]~71_combout ;
wire \rdata_comb[8]~72_combout ;
wire \avl_rddata_local[13]~11_combout ;
wire \avl_rddata_local[13]~10_combout ;
wire \rdata_comb[8]~73_combout ;
wire \csr_flash_cmd_rd_data_0_data[9]~q ;
wire \rdata_comb[9]~74_combout ;
wire \csr_flash_cmd_rd_data_1_data[9]~q ;
wire \rdata_comb[9]~75_combout ;
wire \csr_control_data[9]~q ;
wire \rdata_comb[9]~76_combout ;
wire \csr_flash_cmd_setting_data[9]~q ;
wire \rdata_comb[9]~77_combout ;
wire \rdata_comb[9]~78_combout ;
wire \rdata_comb[9]~79_combout ;
wire \rdata_comb[9]~80_combout ;
wire \csr_flash_cmd_rd_data_0_data[10]~q ;
wire \csr_op_protocol_data[10]~q ;
wire \rdata_comb[10]~81_combout ;
wire \csr_flash_cmd_rd_data_1_data[10]~q ;
wire \rdata_comb[10]~82_combout ;
wire \csr_control_data[10]~q ;
wire \rdata_comb[10]~83_combout ;
wire \csr_flash_cmd_setting_data[10]~q ;
wire \rdata_comb[10]~84_combout ;
wire \rdata_comb[10]~85_combout ;
wire \rdata_comb[10]~86_combout ;
wire \rdata_comb[10]~87_combout ;
wire \csr_flash_cmd_rd_data_0_data[11]~q ;
wire \csr_op_protocol_data[11]~q ;
wire \rdata_comb[11]~88_combout ;
wire \csr_flash_cmd_rd_data_1_data[11]~q ;
wire \rdata_comb[11]~89_combout ;
wire \csr_control_data[11]~q ;
wire \rdata_comb[11]~90_combout ;
wire \csr_flash_cmd_setting_data[11]~2_combout ;
wire \csr_flash_cmd_setting_data[11]~q ;
wire \rdata_comb[11]~91_combout ;
wire \rdata_comb[11]~92_combout ;
wire \rdata_comb[11]~93_combout ;
wire \rdata_comb[11]~94_combout ;
wire \csr_flash_cmd_rd_data_0_data[12]~q ;
wire \rdata_comb[12]~95_combout ;
wire \csr_flash_cmd_rd_data_1_data[12]~q ;
wire \rdata_comb[12]~96_combout ;
wire \csr_control_data[12]~q ;
wire \rdata_comb[12]~97_combout ;
wire \csr_flash_cmd_setting_data[12]~3_combout ;
wire \csr_flash_cmd_setting_data[12]~q ;
wire \rdata_comb[12]~98_combout ;
wire \rdata_comb[12]~99_combout ;
wire \rdata_comb[12]~100_combout ;
wire \rdata_comb[12]~101_combout ;
wire \csr_flash_cmd_rd_data_0_data[13]~q ;
wire \wr_csr_rd_inst~combout ;
wire \csr_rd_inst_data[13]~q ;
wire \rdata_comb[13]~102_combout ;
wire \csr_flash_cmd_rd_data_1_data[13]~q ;
wire \rdata_comb[13]~103_combout ;
wire \csr_control_data[13]~q ;
wire \rdata_comb[13]~104_combout ;
wire \csr_flash_cmd_setting_data[13]~q ;
wire \rdata_comb[13]~105_combout ;
wire \rdata_comb[13]~106_combout ;
wire \rdata_comb[13]~107_combout ;
wire \rdata_comb[13]~108_combout ;
wire \csr_flash_cmd_rd_data_0_data[14]~q ;
wire \csr_rd_inst_data[14]~q ;
wire \csr_op_protocol_data[14]~q ;
wire \rdata_comb[14]~109_combout ;
wire \csr_flash_cmd_rd_data_1_data[14]~q ;
wire \rdata_comb[14]~110_combout ;
wire \csr_control_data[14]~q ;
wire \rdata_comb[14]~111_combout ;
wire \csr_flash_cmd_setting_data[14]~q ;
wire \rdata_comb[14]~112_combout ;
wire \rdata_comb[14]~113_combout ;
wire \rdata_comb[14]~114_combout ;
wire \rdata_comb[14]~115_combout ;
wire \csr_flash_cmd_rd_data_0_data[15]~q ;
wire \csr_rd_inst_data[15]~q ;
wire \csr_op_protocol_data[15]~q ;
wire \rdata_comb[15]~116_combout ;
wire \csr_flash_cmd_rd_data_1_data[15]~q ;
wire \rdata_comb[15]~117_combout ;
wire \csr_control_data[15]~q ;
wire \rdata_comb[15]~118_combout ;
wire \csr_flash_cmd_setting_data[15]~q ;
wire \rdata_comb[15]~119_combout ;
wire \rdata_comb[15]~120_combout ;
wire \rdata_comb[15]~121_combout ;
wire \rdata_comb[15]~122_combout ;
wire \csr_flash_cmd_rd_data_0_data[16]~q ;
wire \csr_rd_inst_data[16]~q ;
wire \rdata_comb[16]~123_combout ;
wire \csr_flash_cmd_rd_data_1_data[16]~q ;
wire \rdata_comb[16]~124_combout ;
wire \csr_control_data[16]~q ;
wire \rdata_comb[16]~125_combout ;
wire \csr_flash_cmd_setting_data[16]~q ;
wire \wr_csr_wr_inst~combout ;
wire \csr_wr_inst_data[16]~q ;
wire \rdata_comb[16]~126_combout ;
wire \rdata_comb[16]~127_combout ;
wire \rdata_comb[16]~128_combout ;
wire \rdata_comb[16]~129_combout ;
wire \csr_flash_cmd_rd_data_0_data[17]~q ;
wire \csr_rd_inst_data[17]~q ;
wire \rdata_comb[17]~130_combout ;
wire \csr_flash_cmd_rd_data_1_data[17]~q ;
wire \rdata_comb[17]~131_combout ;
wire \csr_control_data[17]~q ;
wire \rdata_comb[17]~132_combout ;
wire \csr_flash_cmd_setting_data[17]~q ;
wire \csr_wr_inst_data[17]~q ;
wire \rdata_comb[17]~133_combout ;
wire \rdata_comb[17]~134_combout ;
wire \rdata_comb[17]~135_combout ;
wire \rdata_comb[17]~136_combout ;
wire \csr_rd_inst_data[18]~q ;
wire \csr_flash_cmd_rd_data_0_data[18]~q ;
wire \csr_op_protocol_data[18]~q ;
wire \rdata_comb[18]~137_combout ;
wire \csr_flash_cmd_rd_data_1_data[18]~q ;
wire \rdata_comb[18]~138_combout ;
wire \csr_control_data[18]~q ;
wire \rdata_comb[18]~139_combout ;
wire \csr_flash_cmd_setting_data[18]~q ;
wire \csr_wr_inst_data[18]~q ;
wire \rdata_comb[18]~140_combout ;
wire \rdata_comb[18]~141_combout ;
wire \rdata_comb[18]~142_combout ;
wire \rdata_comb[18]~143_combout ;
wire \csr_rd_inst_data[19]~q ;
wire \csr_flash_cmd_rd_data_0_data[19]~q ;
wire \csr_op_protocol_data[19]~q ;
wire \rdata_comb[19]~144_combout ;
wire \csr_flash_cmd_rd_data_1_data[19]~q ;
wire \rdata_comb[19]~145_combout ;
wire \csr_control_data[19]~q ;
wire \rdata_comb[19]~146_combout ;
wire \csr_flash_cmd_setting_data[19]~q ;
wire \csr_wr_inst_data[19]~q ;
wire \rdata_comb[19]~147_combout ;
wire \rdata_comb[19]~148_combout ;
wire \rdata_comb[19]~149_combout ;
wire \rdata_comb[19]~150_combout ;
wire \csr_rd_inst_data[20]~q ;
wire \csr_flash_cmd_rd_data_0_data[20]~q ;
wire \csr_op_protocol_data[20]~q ;
wire \rdata_comb[20]~151_combout ;
wire \csr_flash_cmd_rd_data_1_data[20]~q ;
wire \rdata_comb[20]~152_combout ;
wire \csr_control_data[20]~q ;
wire \rdata_comb[20]~153_combout ;
wire \csr_flash_cmd_setting_data[20]~q ;
wire \csr_wr_inst_data[20]~q ;
wire \rdata_comb[20]~154_combout ;
wire \rdata_comb[20]~155_combout ;
wire \rdata_comb[20]~156_combout ;
wire \rdata_comb[20]~157_combout ;
wire \csr_rd_inst_data[21]~q ;
wire \csr_flash_cmd_rd_data_0_data[21]~q ;
wire \csr_op_protocol_data[21]~q ;
wire \rdata_comb[21]~158_combout ;
wire \csr_flash_cmd_rd_data_1_data[21]~q ;
wire \rdata_comb[21]~159_combout ;
wire \csr_control_data[21]~q ;
wire \rdata_comb[21]~160_combout ;
wire \csr_flash_cmd_setting_data[21]~q ;
wire \csr_wr_inst_data[21]~q ;
wire \rdata_comb[21]~161_combout ;
wire \rdata_comb[21]~162_combout ;
wire \rdata_comb[21]~163_combout ;
wire \rdata_comb[21]~164_combout ;
wire \csr_rd_inst_data[22]~q ;
wire \csr_flash_cmd_rd_data_0_data[22]~q ;
wire \csr_op_protocol_data[22]~q ;
wire \rdata_comb[22]~165_combout ;
wire \csr_flash_cmd_rd_data_1_data[22]~q ;
wire \rdata_comb[22]~166_combout ;
wire \csr_control_data[22]~q ;
wire \rdata_comb[22]~167_combout ;
wire \csr_flash_cmd_setting_data[22]~q ;
wire \csr_wr_inst_data[22]~q ;
wire \rdata_comb[22]~168_combout ;
wire \rdata_comb[22]~169_combout ;
wire \rdata_comb[22]~170_combout ;
wire \rdata_comb[22]~171_combout ;
wire \csr_rd_inst_data[23]~q ;
wire \csr_flash_cmd_rd_data_0_data[23]~q ;
wire \csr_op_protocol_data[23]~q ;
wire \rdata_comb[23]~172_combout ;
wire \csr_flash_cmd_rd_data_1_data[23]~q ;
wire \rdata_comb[23]~173_combout ;
wire \csr_control_data[23]~q ;
wire \rdata_comb[23]~174_combout ;
wire \csr_flash_cmd_setting_data[23]~q ;
wire \csr_wr_inst_data[23]~q ;
wire \rdata_comb[23]~175_combout ;
wire \rdata_comb[23]~176_combout ;
wire \rdata_comb[23]~177_combout ;
wire \rdata_comb[23]~178_combout ;
wire \csr_rd_inst_data[24]~q ;
wire \csr_flash_cmd_rd_data_0_data[24]~q ;
wire \csr_op_protocol_data[24]~q ;
wire \rdata_comb[24]~179_combout ;
wire \csr_flash_cmd_rd_data_1_data[24]~q ;
wire \rdata_comb[24]~180_combout ;
wire \csr_control_data[24]~q ;
wire \rdata_comb[24]~181_combout ;
wire \csr_flash_cmd_setting_data[24]~q ;
wire \csr_wr_inst_data[24]~q ;
wire \rdata_comb[24]~182_combout ;
wire \rdata_comb[24]~183_combout ;
wire \rdata_comb[24]~184_combout ;
wire \rdata_comb[24]~185_combout ;
wire \csr_rd_inst_data[25]~q ;
wire \csr_flash_cmd_rd_data_0_data[25]~q ;
wire \csr_op_protocol_data[25]~q ;
wire \rdata_comb[25]~186_combout ;
wire \csr_flash_cmd_rd_data_1_data[25]~q ;
wire \rdata_comb[25]~187_combout ;
wire \csr_control_data[25]~q ;
wire \rdata_comb[25]~188_combout ;
wire \csr_flash_cmd_setting_data[25]~q ;
wire \csr_wr_inst_data[25]~q ;
wire \rdata_comb[25]~189_combout ;
wire \rdata_comb[25]~190_combout ;
wire \rdata_comb[25]~191_combout ;
wire \rdata_comb[25]~192_combout ;
wire \csr_rd_inst_data[26]~q ;
wire \csr_flash_cmd_rd_data_0_data[26]~q ;
wire \csr_op_protocol_data[26]~q ;
wire \rdata_comb[26]~193_combout ;
wire \csr_flash_cmd_rd_data_1_data[26]~q ;
wire \rdata_comb[26]~194_combout ;
wire \csr_control_data[26]~q ;
wire \rdata_comb[26]~195_combout ;
wire \csr_flash_cmd_setting_data[26]~q ;
wire \csr_wr_inst_data[26]~q ;
wire \rdata_comb[26]~196_combout ;
wire \rdata_comb[26]~197_combout ;
wire \rdata_comb[26]~198_combout ;
wire \rdata_comb[26]~199_combout ;
wire \csr_rd_inst_data[27]~q ;
wire \csr_flash_cmd_rd_data_0_data[27]~q ;
wire \csr_op_protocol_data[27]~q ;
wire \rdata_comb[27]~200_combout ;
wire \csr_flash_cmd_rd_data_1_data[27]~q ;
wire \rdata_comb[27]~201_combout ;
wire \csr_control_data[27]~q ;
wire \rdata_comb[27]~202_combout ;
wire \csr_flash_cmd_setting_data[27]~q ;
wire \csr_wr_inst_data[27]~q ;
wire \rdata_comb[27]~203_combout ;
wire \rdata_comb[27]~204_combout ;
wire \rdata_comb[27]~205_combout ;
wire \rdata_comb[27]~206_combout ;
wire \csr_rd_inst_data[28]~q ;
wire \csr_flash_cmd_rd_data_0_data[28]~q ;
wire \csr_op_protocol_data[28]~q ;
wire \rdata_comb[28]~207_combout ;
wire \csr_flash_cmd_rd_data_1_data[28]~q ;
wire \rdata_comb[28]~208_combout ;
wire \csr_control_data[28]~q ;
wire \rdata_comb[28]~209_combout ;
wire \csr_flash_cmd_setting_data[28]~q ;
wire \csr_wr_inst_data[28]~q ;
wire \rdata_comb[28]~210_combout ;
wire \rdata_comb[28]~211_combout ;
wire \rdata_comb[28]~212_combout ;
wire \rdata_comb[28]~213_combout ;
wire \csr_rd_inst_data[29]~q ;
wire \csr_flash_cmd_rd_data_0_data[29]~q ;
wire \csr_op_protocol_data[29]~q ;
wire \rdata_comb[29]~214_combout ;
wire \csr_flash_cmd_rd_data_1_data[29]~q ;
wire \rdata_comb[29]~215_combout ;
wire \csr_control_data[29]~q ;
wire \rdata_comb[29]~216_combout ;
wire \csr_flash_cmd_setting_data[29]~q ;
wire \csr_wr_inst_data[29]~q ;
wire \rdata_comb[29]~217_combout ;
wire \rdata_comb[29]~218_combout ;
wire \rdata_comb[29]~219_combout ;
wire \rdata_comb[29]~220_combout ;
wire \csr_rd_inst_data[30]~q ;
wire \csr_flash_cmd_rd_data_0_data[30]~q ;
wire \csr_op_protocol_data[30]~q ;
wire \rdata_comb[30]~221_combout ;
wire \csr_flash_cmd_rd_data_1_data[30]~q ;
wire \rdata_comb[30]~222_combout ;
wire \csr_control_data[30]~q ;
wire \rdata_comb[30]~223_combout ;
wire \csr_flash_cmd_setting_data[30]~q ;
wire \csr_wr_inst_data[30]~q ;
wire \rdata_comb[30]~224_combout ;
wire \rdata_comb[30]~225_combout ;
wire \rdata_comb[30]~226_combout ;
wire \rdata_comb[30]~227_combout ;
wire \csr_rd_inst_data[31]~q ;
wire \csr_flash_cmd_rd_data_0_data[31]~q ;
wire \csr_op_protocol_data[31]~q ;
wire \rdata_comb[31]~228_combout ;
wire \csr_flash_cmd_rd_data_1_data[31]~q ;
wire \rdata_comb[31]~229_combout ;
wire \csr_control_data[31]~q ;
wire \rdata_comb[31]~230_combout ;
wire \csr_flash_cmd_setting_data[31]~q ;
wire \csr_wr_inst_data[31]~q ;
wire \rdata_comb[31]~231_combout ;
wire \rdata_comb[31]~232_combout ;
wire \rdata_comb[31]~233_combout ;
wire \rdata_comb[31]~234_combout ;
wire \Selector32~0_combout ;
wire \wr_csr_flash_cmd_control~0_combout ;
wire \wr_csr_flash_cmd_control~1_combout ;
wire \wr_csr_flash_cmd_control~2_combout ;
wire \wr_csr_flash_cmd_control~3_combout ;
wire \wr_csr_flash_cmd_control~4_combout ;
wire \wr_csr_flash_cmd_control~5_combout ;
wire \wr_csr_flash_cmd_control~6_combout ;
wire \wr_csr_flash_cmd_control~7_combout ;
wire \wr_csr_flash_cmd_control~8_combout ;
wire \wr_csr_flash_cmd_control~9_combout ;
wire \wr_csr_flash_cmd_control~10_combout ;
wire \wr_csr_flash_cmd_control~11_combout ;
wire \flash_operation_reg~q ;
wire \Selector32~1_combout ;
wire \avl_rddatavalid_local~0_combout ;
wire \csr_rd_inst_data[0]~0_combout ;
wire \wr_csr_flash_cmd_wr_data_0~combout ;
wire \wr_csr_flash_cmd_addr~combout ;
wire \wr_csr_flash_cmd_wr_data_1~combout ;
wire \wr_csr_delay_setting~combout ;
wire \csr_clk_baud_rate_data[4]~2_combout ;
wire \csr_clk_baud_rate_data[4]~4_combout ;
wire \csr_clk_baud_rate_data[4]~3_combout ;
wire \csr_control_data[0]~0_combout ;
wire \wr_csr_rd_capturing~combout ;
wire \csr_wr_inst_data[1]~0_combout ;
wire \csr_rd_inst_data[1]~1_combout ;
wire \csr_clk_baud_rate_data[4]~5_combout ;
wire \csr_wr_inst_data[12]~1_combout ;
wire \csr_wr_inst_data[13]~2_combout ;
wire \csr_wr_inst_data[14]~3_combout ;
wire \Selector36~0_combout ;
wire \Selector36~1_combout ;
wire \Selector33~0_combout ;
wire \Selector35~0_combout ;
wire \Equal16~0_combout ;
wire \has_data_in~0_combout ;
wire \LessThan0~0_combout ;
wire \has_data_out~0_combout ;
wire \numb_data[0]~0_combout ;
wire \Equal13~0_combout ;
wire \Equal14~0_combout ;
wire \opcode[0]~0_combout ;
wire \opcode[2]~1_combout ;
wire \Equal15~0_combout ;
wire \Equal15~1_combout ;


dffeas \avl_rddata_local[0] (
	.clk(clk),
	.d(\rdata_comb[0]~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_0),
	.prn(vcc));
defparam \avl_rddata_local[0] .is_wysiwyg = "true";
defparam \avl_rddata_local[0] .power_up = "low";

dffeas \avl_rddata_local[1] (
	.clk(clk),
	.d(\rdata_comb[1]~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_1),
	.prn(vcc));
defparam \avl_rddata_local[1] .is_wysiwyg = "true";
defparam \avl_rddata_local[1] .power_up = "low";

dffeas \avl_rddata_local[2] (
	.clk(clk),
	.d(\rdata_comb[2]~29_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_2),
	.prn(vcc));
defparam \avl_rddata_local[2] .is_wysiwyg = "true";
defparam \avl_rddata_local[2] .power_up = "low";

dffeas \avl_rddata_local[3] (
	.clk(clk),
	.d(\rdata_comb[3]~38_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_3),
	.prn(vcc));
defparam \avl_rddata_local[3] .is_wysiwyg = "true";
defparam \avl_rddata_local[3] .power_up = "low";

dffeas \avl_rddata_local[4] (
	.clk(clk),
	.d(\rdata_comb[4]~235_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_4),
	.prn(vcc));
defparam \avl_rddata_local[4] .is_wysiwyg = "true";
defparam \avl_rddata_local[4] .power_up = "low";

dffeas \avl_rddata_local[5] (
	.clk(clk),
	.d(\rdata_comb[5]~48_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_5),
	.prn(vcc));
defparam \avl_rddata_local[5] .is_wysiwyg = "true";
defparam \avl_rddata_local[5] .power_up = "low";

dffeas \avl_rddata_local[6] (
	.clk(clk),
	.d(\rdata_comb[6]~57_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_6),
	.prn(vcc));
defparam \avl_rddata_local[6] .is_wysiwyg = "true";
defparam \avl_rddata_local[6] .power_up = "low";

dffeas \avl_rddata_local[7] (
	.clk(clk),
	.d(\rdata_comb[7]~66_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_7),
	.prn(vcc));
defparam \avl_rddata_local[7] .is_wysiwyg = "true";
defparam \avl_rddata_local[7] .power_up = "low";

dffeas \avl_rddata_local[8] (
	.clk(clk),
	.d(\rdata_comb[8]~73_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_8),
	.prn(vcc));
defparam \avl_rddata_local[8] .is_wysiwyg = "true";
defparam \avl_rddata_local[8] .power_up = "low";

dffeas \avl_rddata_local[9] (
	.clk(clk),
	.d(\rdata_comb[9]~80_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_9),
	.prn(vcc));
defparam \avl_rddata_local[9] .is_wysiwyg = "true";
defparam \avl_rddata_local[9] .power_up = "low";

dffeas \avl_rddata_local[10] (
	.clk(clk),
	.d(\rdata_comb[10]~87_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_10),
	.prn(vcc));
defparam \avl_rddata_local[10] .is_wysiwyg = "true";
defparam \avl_rddata_local[10] .power_up = "low";

dffeas \avl_rddata_local[11] (
	.clk(clk),
	.d(\rdata_comb[11]~94_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_11),
	.prn(vcc));
defparam \avl_rddata_local[11] .is_wysiwyg = "true";
defparam \avl_rddata_local[11] .power_up = "low";

dffeas \avl_rddata_local[12] (
	.clk(clk),
	.d(\rdata_comb[12]~101_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_12),
	.prn(vcc));
defparam \avl_rddata_local[12] .is_wysiwyg = "true";
defparam \avl_rddata_local[12] .power_up = "low";

dffeas \avl_rddata_local[13] (
	.clk(clk),
	.d(\rdata_comb[13]~108_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_13),
	.prn(vcc));
defparam \avl_rddata_local[13] .is_wysiwyg = "true";
defparam \avl_rddata_local[13] .power_up = "low";

dffeas \avl_rddata_local[14] (
	.clk(clk),
	.d(\rdata_comb[14]~115_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_14),
	.prn(vcc));
defparam \avl_rddata_local[14] .is_wysiwyg = "true";
defparam \avl_rddata_local[14] .power_up = "low";

dffeas \avl_rddata_local[15] (
	.clk(clk),
	.d(\rdata_comb[15]~122_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_15),
	.prn(vcc));
defparam \avl_rddata_local[15] .is_wysiwyg = "true";
defparam \avl_rddata_local[15] .power_up = "low";

dffeas \avl_rddata_local[16] (
	.clk(clk),
	.d(\rdata_comb[16]~129_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_16),
	.prn(vcc));
defparam \avl_rddata_local[16] .is_wysiwyg = "true";
defparam \avl_rddata_local[16] .power_up = "low";

dffeas \avl_rddata_local[17] (
	.clk(clk),
	.d(\rdata_comb[17]~136_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_17),
	.prn(vcc));
defparam \avl_rddata_local[17] .is_wysiwyg = "true";
defparam \avl_rddata_local[17] .power_up = "low";

dffeas \avl_rddata_local[18] (
	.clk(clk),
	.d(\rdata_comb[18]~143_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_18),
	.prn(vcc));
defparam \avl_rddata_local[18] .is_wysiwyg = "true";
defparam \avl_rddata_local[18] .power_up = "low";

dffeas \avl_rddata_local[19] (
	.clk(clk),
	.d(\rdata_comb[19]~150_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_19),
	.prn(vcc));
defparam \avl_rddata_local[19] .is_wysiwyg = "true";
defparam \avl_rddata_local[19] .power_up = "low";

dffeas \avl_rddata_local[20] (
	.clk(clk),
	.d(\rdata_comb[20]~157_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_20),
	.prn(vcc));
defparam \avl_rddata_local[20] .is_wysiwyg = "true";
defparam \avl_rddata_local[20] .power_up = "low";

dffeas \avl_rddata_local[21] (
	.clk(clk),
	.d(\rdata_comb[21]~164_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_21),
	.prn(vcc));
defparam \avl_rddata_local[21] .is_wysiwyg = "true";
defparam \avl_rddata_local[21] .power_up = "low";

dffeas \avl_rddata_local[22] (
	.clk(clk),
	.d(\rdata_comb[22]~171_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_22),
	.prn(vcc));
defparam \avl_rddata_local[22] .is_wysiwyg = "true";
defparam \avl_rddata_local[22] .power_up = "low";

dffeas \avl_rddata_local[23] (
	.clk(clk),
	.d(\rdata_comb[23]~178_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_23),
	.prn(vcc));
defparam \avl_rddata_local[23] .is_wysiwyg = "true";
defparam \avl_rddata_local[23] .power_up = "low";

dffeas \avl_rddata_local[24] (
	.clk(clk),
	.d(\rdata_comb[24]~185_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_24),
	.prn(vcc));
defparam \avl_rddata_local[24] .is_wysiwyg = "true";
defparam \avl_rddata_local[24] .power_up = "low";

dffeas \avl_rddata_local[25] (
	.clk(clk),
	.d(\rdata_comb[25]~192_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_25),
	.prn(vcc));
defparam \avl_rddata_local[25] .is_wysiwyg = "true";
defparam \avl_rddata_local[25] .power_up = "low";

dffeas \avl_rddata_local[26] (
	.clk(clk),
	.d(\rdata_comb[26]~199_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_26),
	.prn(vcc));
defparam \avl_rddata_local[26] .is_wysiwyg = "true";
defparam \avl_rddata_local[26] .power_up = "low";

dffeas \avl_rddata_local[27] (
	.clk(clk),
	.d(\rdata_comb[27]~206_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_27),
	.prn(vcc));
defparam \avl_rddata_local[27] .is_wysiwyg = "true";
defparam \avl_rddata_local[27] .power_up = "low";

dffeas \avl_rddata_local[28] (
	.clk(clk),
	.d(\rdata_comb[28]~213_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_28),
	.prn(vcc));
defparam \avl_rddata_local[28] .is_wysiwyg = "true";
defparam \avl_rddata_local[28] .power_up = "low";

dffeas \avl_rddata_local[29] (
	.clk(clk),
	.d(\rdata_comb[29]~220_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_29),
	.prn(vcc));
defparam \avl_rddata_local[29] .is_wysiwyg = "true";
defparam \avl_rddata_local[29] .power_up = "low";

dffeas \avl_rddata_local[30] (
	.clk(clk),
	.d(\rdata_comb[30]~227_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_30),
	.prn(vcc));
defparam \avl_rddata_local[30] .is_wysiwyg = "true";
defparam \avl_rddata_local[30] .power_up = "low";

dffeas \avl_rddata_local[31] (
	.clk(clk),
	.d(\rdata_comb[31]~234_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddata_local_31),
	.prn(vcc));
defparam \avl_rddata_local[31] .is_wysiwyg = "true";
defparam \avl_rddata_local[31] .power_up = "low";

dffeas \state.ST_IDLE (
	.clk(clk),
	.d(\Selector32~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stateST_IDLE),
	.prn(vcc));
defparam \state.ST_IDLE .is_wysiwyg = "true";
defparam \state.ST_IDLE .power_up = "low";

cycloneive_lcell_comb csr_waitrequest(
	.dataa(\flash_operation_reg~q ),
	.datab(stateST_IDLE),
	.datac(gnd),
	.datad(hold_waitrequest),
	.cin(gnd),
	.combout(csr_waitrequest1),
	.cout());
defparam csr_waitrequest.lut_mask = 16'hEEFF;
defparam csr_waitrequest.sum_lutc_input = "datac";

dffeas avl_rddatavalid_local(
	.clk(clk),
	.d(\avl_rddatavalid_local~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(avl_rddatavalid_local1),
	.prn(vcc));
defparam avl_rddatavalid_local.is_wysiwyg = "true";
defparam avl_rddatavalid_local.power_up = "low";

dffeas \csr_wr_inst_data[0] (
	.clk(clk),
	.d(csr_wrdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(csr_wr_inst_data_0),
	.prn(vcc));
defparam \csr_wr_inst_data[0] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[0] .power_up = "low";

dffeas \csr_rd_inst_data[0] (
	.clk(clk),
	.d(\csr_rd_inst_data[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(csr_rd_inst_data_0),
	.prn(vcc));
defparam \csr_rd_inst_data[0] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[0] .power_up = "low";

dffeas \csr_op_protocol_data[0] (
	.clk(clk),
	.d(csr_wrdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(csr_op_protocol_data_0),
	.prn(vcc));
defparam \csr_op_protocol_data[0] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[0] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[0] (
	.clk(clk),
	.d(csr_wrdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_0),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[0] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[0] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[0] (
	.clk(clk),
	.d(csr_wrdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_0),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[0] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[0] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[0] (
	.clk(clk),
	.d(csr_wrdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_0),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[0] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[0] .power_up = "low";

dffeas \csr_delay_setting_data[0] (
	.clk(clk),
	.d(csr_wrdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_delay_setting~combout ),
	.q(csr_delay_setting_data_0),
	.prn(vcc));
defparam \csr_delay_setting_data[0] .is_wysiwyg = "true";
defparam \csr_delay_setting_data[0] .power_up = "low";

dffeas \csr_clk_baud_rate_data[0] (
	.clk(clk),
	.d(csr_wrdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_clk_baud_rate_data[4]~3_combout ),
	.q(csr_clk_baud_rate_data_0),
	.prn(vcc));
defparam \csr_clk_baud_rate_data[0] .is_wysiwyg = "true";
defparam \csr_clk_baud_rate_data[0] .power_up = "low";

dffeas \csr_control_data[0] (
	.clk(clk),
	.d(\csr_control_data[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(csr_control_data_0),
	.prn(vcc));
defparam \csr_control_data[0] .is_wysiwyg = "true";
defparam \csr_control_data[0] .power_up = "low";

dffeas \csr_rd_capturing_data[0] (
	.clk(clk),
	.d(csr_wrdata[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_capturing~combout ),
	.q(csr_rd_capturing_data_0),
	.prn(vcc));
defparam \csr_rd_capturing_data[0] .is_wysiwyg = "true";
defparam \csr_rd_capturing_data[0] .power_up = "low";

dffeas \csr_wr_inst_data[1] (
	.clk(clk),
	.d(\csr_wr_inst_data[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(csr_wr_inst_data_1),
	.prn(vcc));
defparam \csr_wr_inst_data[1] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[1] .power_up = "low";

dffeas \csr_rd_inst_data[1] (
	.clk(clk),
	.d(\csr_rd_inst_data[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(csr_rd_inst_data_1),
	.prn(vcc));
defparam \csr_rd_inst_data[1] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[1] .power_up = "low";

dffeas \csr_op_protocol_data[1] (
	.clk(clk),
	.d(csr_wrdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(csr_op_protocol_data_1),
	.prn(vcc));
defparam \csr_op_protocol_data[1] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[1] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[1] (
	.clk(clk),
	.d(csr_wrdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_1),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[1] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[1] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[1] (
	.clk(clk),
	.d(csr_wrdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_1),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[1] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[1] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[1] (
	.clk(clk),
	.d(csr_wrdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_1),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[1] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[1] .power_up = "low";

dffeas \csr_delay_setting_data[1] (
	.clk(clk),
	.d(csr_wrdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_delay_setting~combout ),
	.q(csr_delay_setting_data_1),
	.prn(vcc));
defparam \csr_delay_setting_data[1] .is_wysiwyg = "true";
defparam \csr_delay_setting_data[1] .power_up = "low";

dffeas \csr_clk_baud_rate_data[1] (
	.clk(clk),
	.d(csr_wrdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_clk_baud_rate_data[4]~3_combout ),
	.q(csr_clk_baud_rate_data_1),
	.prn(vcc));
defparam \csr_clk_baud_rate_data[1] .is_wysiwyg = "true";
defparam \csr_clk_baud_rate_data[1] .power_up = "low";

dffeas \csr_rd_capturing_data[1] (
	.clk(clk),
	.d(csr_wrdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_capturing~combout ),
	.q(csr_rd_capturing_data_1),
	.prn(vcc));
defparam \csr_rd_capturing_data[1] .is_wysiwyg = "true";
defparam \csr_rd_capturing_data[1] .power_up = "low";

dffeas \csr_wr_inst_data[2] (
	.clk(clk),
	.d(csr_wrdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(csr_wr_inst_data_2),
	.prn(vcc));
defparam \csr_wr_inst_data[2] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[2] .power_up = "low";

dffeas \csr_rd_inst_data[2] (
	.clk(clk),
	.d(csr_wrdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(csr_rd_inst_data_2),
	.prn(vcc));
defparam \csr_rd_inst_data[2] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[2] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[2] (
	.clk(clk),
	.d(csr_wrdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_2),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[2] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[2] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[2] (
	.clk(clk),
	.d(csr_wrdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_2),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[2] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[2] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[2] (
	.clk(clk),
	.d(csr_wrdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_2),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[2] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[2] .power_up = "low";

dffeas \csr_delay_setting_data[2] (
	.clk(clk),
	.d(csr_wrdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_delay_setting~combout ),
	.q(csr_delay_setting_data_2),
	.prn(vcc));
defparam \csr_delay_setting_data[2] .is_wysiwyg = "true";
defparam \csr_delay_setting_data[2] .power_up = "low";

dffeas \csr_clk_baud_rate_data[2] (
	.clk(clk),
	.d(csr_wrdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_clk_baud_rate_data[4]~3_combout ),
	.q(csr_clk_baud_rate_data_2),
	.prn(vcc));
defparam \csr_clk_baud_rate_data[2] .is_wysiwyg = "true";
defparam \csr_clk_baud_rate_data[2] .power_up = "low";

dffeas \csr_rd_capturing_data[2] (
	.clk(clk),
	.d(csr_wrdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_capturing~combout ),
	.q(csr_rd_capturing_data_2),
	.prn(vcc));
defparam \csr_rd_capturing_data[2] .is_wysiwyg = "true";
defparam \csr_rd_capturing_data[2] .power_up = "low";

dffeas \csr_wr_inst_data[3] (
	.clk(clk),
	.d(csr_wrdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(csr_wr_inst_data_3),
	.prn(vcc));
defparam \csr_wr_inst_data[3] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[3] .power_up = "low";

dffeas \csr_rd_inst_data[3] (
	.clk(clk),
	.d(csr_wrdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(csr_rd_inst_data_3),
	.prn(vcc));
defparam \csr_rd_inst_data[3] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[3] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[3] (
	.clk(clk),
	.d(csr_wrdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_3),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[3] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[3] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[3] (
	.clk(clk),
	.d(csr_wrdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_3),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[3] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[3] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[3] (
	.clk(clk),
	.d(csr_wrdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_3),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[3] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[3] .power_up = "low";

dffeas \csr_delay_setting_data[3] (
	.clk(clk),
	.d(csr_wrdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_delay_setting~combout ),
	.q(csr_delay_setting_data_3),
	.prn(vcc));
defparam \csr_delay_setting_data[3] .is_wysiwyg = "true";
defparam \csr_delay_setting_data[3] .power_up = "low";

dffeas \csr_clk_baud_rate_data[3] (
	.clk(clk),
	.d(csr_wrdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_clk_baud_rate_data[4]~3_combout ),
	.q(csr_clk_baud_rate_data_3),
	.prn(vcc));
defparam \csr_clk_baud_rate_data[3] .is_wysiwyg = "true";
defparam \csr_clk_baud_rate_data[3] .power_up = "low";

dffeas \csr_rd_capturing_data[3] (
	.clk(clk),
	.d(csr_wrdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_capturing~combout ),
	.q(csr_rd_capturing_data_3),
	.prn(vcc));
defparam \csr_rd_capturing_data[3] .is_wysiwyg = "true";
defparam \csr_rd_capturing_data[3] .power_up = "low";

dffeas \csr_wr_inst_data[4] (
	.clk(clk),
	.d(csr_wrdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(csr_wr_inst_data_4),
	.prn(vcc));
defparam \csr_wr_inst_data[4] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[4] .power_up = "low";

dffeas \csr_delay_setting_data[4] (
	.clk(clk),
	.d(csr_wrdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_delay_setting~combout ),
	.q(csr_delay_setting_data_4),
	.prn(vcc));
defparam \csr_delay_setting_data[4] .is_wysiwyg = "true";
defparam \csr_delay_setting_data[4] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[4] (
	.clk(clk),
	.d(csr_wrdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_4),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[4] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[4] .power_up = "low";

dffeas \csr_op_protocol_data[4] (
	.clk(clk),
	.d(csr_wrdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(csr_op_protocol_data_4),
	.prn(vcc));
defparam \csr_op_protocol_data[4] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[4] .power_up = "low";

dffeas \csr_clk_baud_rate_data[4] (
	.clk(clk),
	.d(\csr_clk_baud_rate_data[4]~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_clk_baud_rate_data[4]~3_combout ),
	.q(csr_clk_baud_rate_data_4),
	.prn(vcc));
defparam \csr_clk_baud_rate_data[4] .is_wysiwyg = "true";
defparam \csr_clk_baud_rate_data[4] .power_up = "low";

dffeas \csr_control_data[4] (
	.clk(clk),
	.d(csr_wrdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(csr_control_data_4),
	.prn(vcc));
defparam \csr_control_data[4] .is_wysiwyg = "true";
defparam \csr_control_data[4] .power_up = "low";

dffeas \csr_rd_inst_data[4] (
	.clk(clk),
	.d(csr_wrdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(csr_rd_inst_data_4),
	.prn(vcc));
defparam \csr_rd_inst_data[4] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[4] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[4] (
	.clk(clk),
	.d(csr_wrdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_4),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[4] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[4] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[4] (
	.clk(clk),
	.d(csr_wrdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_4),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[4] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[4] .power_up = "low";

dffeas \csr_delay_setting_data[5] (
	.clk(clk),
	.d(csr_wrdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_delay_setting~combout ),
	.q(csr_delay_setting_data_5),
	.prn(vcc));
defparam \csr_delay_setting_data[5] .is_wysiwyg = "true";
defparam \csr_delay_setting_data[5] .power_up = "low";

dffeas \csr_wr_inst_data[5] (
	.clk(clk),
	.d(csr_wrdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(csr_wr_inst_data_5),
	.prn(vcc));
defparam \csr_wr_inst_data[5] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[5] .power_up = "low";

dffeas \csr_rd_inst_data[5] (
	.clk(clk),
	.d(csr_wrdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(csr_rd_inst_data_5),
	.prn(vcc));
defparam \csr_rd_inst_data[5] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[5] .power_up = "low";

dffeas \csr_op_protocol_data[5] (
	.clk(clk),
	.d(csr_wrdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(csr_op_protocol_data_5),
	.prn(vcc));
defparam \csr_op_protocol_data[5] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[5] .power_up = "low";

dffeas \csr_control_data[5] (
	.clk(clk),
	.d(csr_wrdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(csr_control_data_5),
	.prn(vcc));
defparam \csr_control_data[5] .is_wysiwyg = "true";
defparam \csr_control_data[5] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[5] (
	.clk(clk),
	.d(csr_wrdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_5),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[5] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[5] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[5] (
	.clk(clk),
	.d(csr_wrdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_5),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[5] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[5] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[5] (
	.clk(clk),
	.d(csr_wrdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_5),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[5] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[5] .power_up = "low";

dffeas \csr_wr_inst_data[6] (
	.clk(clk),
	.d(csr_wrdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(csr_wr_inst_data_6),
	.prn(vcc));
defparam \csr_wr_inst_data[6] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[6] .power_up = "low";

dffeas \csr_rd_inst_data[6] (
	.clk(clk),
	.d(csr_wrdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(csr_rd_inst_data_6),
	.prn(vcc));
defparam \csr_rd_inst_data[6] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[6] .power_up = "low";

dffeas \csr_delay_setting_data[6] (
	.clk(clk),
	.d(csr_wrdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_delay_setting~combout ),
	.q(csr_delay_setting_data_6),
	.prn(vcc));
defparam \csr_delay_setting_data[6] .is_wysiwyg = "true";
defparam \csr_delay_setting_data[6] .power_up = "low";

dffeas \csr_control_data[6] (
	.clk(clk),
	.d(csr_wrdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(csr_control_data_6),
	.prn(vcc));
defparam \csr_control_data[6] .is_wysiwyg = "true";
defparam \csr_control_data[6] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[6] (
	.clk(clk),
	.d(csr_wrdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_6),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[6] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[6] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[6] (
	.clk(clk),
	.d(csr_wrdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_6),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[6] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[6] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[6] (
	.clk(clk),
	.d(csr_wrdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_6),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[6] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[6] .power_up = "low";

dffeas \csr_delay_setting_data[7] (
	.clk(clk),
	.d(csr_wrdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_delay_setting~combout ),
	.q(csr_delay_setting_data_7),
	.prn(vcc));
defparam \csr_delay_setting_data[7] .is_wysiwyg = "true";
defparam \csr_delay_setting_data[7] .power_up = "low";

dffeas \csr_wr_inst_data[7] (
	.clk(clk),
	.d(csr_wrdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(csr_wr_inst_data_7),
	.prn(vcc));
defparam \csr_wr_inst_data[7] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[7] .power_up = "low";

dffeas \csr_rd_inst_data[7] (
	.clk(clk),
	.d(csr_wrdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(csr_rd_inst_data_7),
	.prn(vcc));
defparam \csr_rd_inst_data[7] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[7] .power_up = "low";

dffeas \csr_control_data[7] (
	.clk(clk),
	.d(csr_wrdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(csr_control_data_7),
	.prn(vcc));
defparam \csr_control_data[7] .is_wysiwyg = "true";
defparam \csr_control_data[7] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[7] (
	.clk(clk),
	.d(csr_wrdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_7),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[7] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[7] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[7] (
	.clk(clk),
	.d(csr_wrdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_7),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[7] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[7] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[7] (
	.clk(clk),
	.d(csr_wrdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_7),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[7] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[7] .power_up = "low";

dffeas \csr_rd_inst_data[8] (
	.clk(clk),
	.d(csr_wrdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(csr_rd_inst_data_8),
	.prn(vcc));
defparam \csr_rd_inst_data[8] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[8] .power_up = "low";

dffeas \csr_op_protocol_data[8] (
	.clk(clk),
	.d(csr_wrdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(csr_op_protocol_data_8),
	.prn(vcc));
defparam \csr_op_protocol_data[8] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[8] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[8] (
	.clk(clk),
	.d(csr_wrdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_8),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[8] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[8] .power_up = "low";

dffeas \csr_control_data[8] (
	.clk(clk),
	.d(csr_wrdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(csr_control_data_8),
	.prn(vcc));
defparam \csr_control_data[8] .is_wysiwyg = "true";
defparam \csr_control_data[8] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[8] (
	.clk(clk),
	.d(csr_wrdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_8),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[8] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[8] .power_up = "low";

dffeas \csr_wr_inst_data[8] (
	.clk(clk),
	.d(csr_wrdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(csr_wr_inst_data_8),
	.prn(vcc));
defparam \csr_wr_inst_data[8] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[8] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[8] (
	.clk(clk),
	.d(csr_wrdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_8),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[8] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[8] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[9] (
	.clk(clk),
	.d(csr_wrdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_9),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[9] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[9] .power_up = "low";

dffeas \csr_rd_inst_data[9] (
	.clk(clk),
	.d(csr_wrdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(csr_rd_inst_data_9),
	.prn(vcc));
defparam \csr_rd_inst_data[9] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[9] .power_up = "low";

dffeas \csr_op_protocol_data[9] (
	.clk(clk),
	.d(csr_wrdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(csr_op_protocol_data_9),
	.prn(vcc));
defparam \csr_op_protocol_data[9] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[9] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[9] (
	.clk(clk),
	.d(csr_wrdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_9),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[9] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[9] .power_up = "low";

dffeas \csr_wr_inst_data[9] (
	.clk(clk),
	.d(csr_wrdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(csr_wr_inst_data_9),
	.prn(vcc));
defparam \csr_wr_inst_data[9] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[9] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[9] (
	.clk(clk),
	.d(csr_wrdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_9),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[9] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[9] .power_up = "low";

dffeas \csr_rd_inst_data[10] (
	.clk(clk),
	.d(csr_wrdata[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(csr_rd_inst_data_10),
	.prn(vcc));
defparam \csr_rd_inst_data[10] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[10] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[10] (
	.clk(clk),
	.d(csr_wrdata[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_10),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[10] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[10] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[10] (
	.clk(clk),
	.d(csr_wrdata[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_10),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[10] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[10] .power_up = "low";

dffeas \csr_wr_inst_data[10] (
	.clk(clk),
	.d(csr_wrdata[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(csr_wr_inst_data_10),
	.prn(vcc));
defparam \csr_wr_inst_data[10] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[10] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[10] (
	.clk(clk),
	.d(csr_wrdata[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_10),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[10] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[10] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[11] (
	.clk(clk),
	.d(csr_wrdata[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_11),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[11] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[11] .power_up = "low";

dffeas \csr_rd_inst_data[11] (
	.clk(clk),
	.d(csr_wrdata[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(csr_rd_inst_data_11),
	.prn(vcc));
defparam \csr_rd_inst_data[11] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[11] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[11] (
	.clk(clk),
	.d(csr_wrdata[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_11),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[11] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[11] .power_up = "low";

dffeas \csr_wr_inst_data[11] (
	.clk(clk),
	.d(csr_wrdata[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(csr_wr_inst_data_11),
	.prn(vcc));
defparam \csr_wr_inst_data[11] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[11] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[11] (
	.clk(clk),
	.d(csr_wrdata[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_11),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[11] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[11] .power_up = "low";

dffeas \csr_rd_inst_data[12] (
	.clk(clk),
	.d(csr_wrdata[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(csr_rd_inst_data_12),
	.prn(vcc));
defparam \csr_rd_inst_data[12] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[12] .power_up = "low";

dffeas \csr_op_protocol_data[12] (
	.clk(clk),
	.d(csr_wrdata[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(csr_op_protocol_data_12),
	.prn(vcc));
defparam \csr_op_protocol_data[12] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[12] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[12] (
	.clk(clk),
	.d(csr_wrdata[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_12),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[12] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[12] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[12] (
	.clk(clk),
	.d(csr_wrdata[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_12),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[12] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[12] .power_up = "low";

dffeas \csr_wr_inst_data[12] (
	.clk(clk),
	.d(\csr_wr_inst_data[12]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(csr_wr_inst_data_12),
	.prn(vcc));
defparam \csr_wr_inst_data[12] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[12] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[12] (
	.clk(clk),
	.d(csr_wrdata[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_12),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[12] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[12] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[13] (
	.clk(clk),
	.d(csr_wrdata[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_13),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[13] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[13] .power_up = "low";

dffeas \csr_op_protocol_data[13] (
	.clk(clk),
	.d(csr_wrdata[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(csr_op_protocol_data_13),
	.prn(vcc));
defparam \csr_op_protocol_data[13] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[13] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[13] (
	.clk(clk),
	.d(csr_wrdata[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_13),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[13] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[13] .power_up = "low";

dffeas \csr_wr_inst_data[13] (
	.clk(clk),
	.d(\csr_wr_inst_data[13]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(csr_wr_inst_data_13),
	.prn(vcc));
defparam \csr_wr_inst_data[13] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[13] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[13] (
	.clk(clk),
	.d(csr_wrdata[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_13),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[13] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[13] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[14] (
	.clk(clk),
	.d(csr_wrdata[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_14),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[14] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[14] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[14] (
	.clk(clk),
	.d(csr_wrdata[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_14),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[14] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[14] .power_up = "low";

dffeas \csr_wr_inst_data[14] (
	.clk(clk),
	.d(\csr_wr_inst_data[14]~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(csr_wr_inst_data_14),
	.prn(vcc));
defparam \csr_wr_inst_data[14] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[14] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[14] (
	.clk(clk),
	.d(csr_wrdata[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_14),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[14] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[14] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[15] (
	.clk(clk),
	.d(csr_wrdata[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_15),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[15] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[15] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[15] (
	.clk(clk),
	.d(csr_wrdata[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_15),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[15] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[15] .power_up = "low";

dffeas \csr_wr_inst_data[15] (
	.clk(clk),
	.d(csr_wrdata[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(csr_wr_inst_data_15),
	.prn(vcc));
defparam \csr_wr_inst_data[15] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[15] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[15] (
	.clk(clk),
	.d(csr_wrdata[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_15),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[15] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[15] .power_up = "low";

dffeas \csr_op_protocol_data[16] (
	.clk(clk),
	.d(csr_wrdata[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(csr_op_protocol_data_16),
	.prn(vcc));
defparam \csr_op_protocol_data[16] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[16] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[16] (
	.clk(clk),
	.d(csr_wrdata[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_16),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[16] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[16] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[16] (
	.clk(clk),
	.d(csr_wrdata[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_16),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[16] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[16] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[16] (
	.clk(clk),
	.d(csr_wrdata[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_16),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[16] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[16] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[17] (
	.clk(clk),
	.d(csr_wrdata[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_17),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[17] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[17] .power_up = "low";

dffeas \csr_op_protocol_data[17] (
	.clk(clk),
	.d(csr_wrdata[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(csr_op_protocol_data_17),
	.prn(vcc));
defparam \csr_op_protocol_data[17] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[17] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[17] (
	.clk(clk),
	.d(csr_wrdata[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_17),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[17] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[17] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[17] (
	.clk(clk),
	.d(csr_wrdata[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_17),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[17] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[17] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[18] (
	.clk(clk),
	.d(csr_wrdata[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_18),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[18] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[18] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[18] (
	.clk(clk),
	.d(csr_wrdata[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_18),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[18] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[18] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[18] (
	.clk(clk),
	.d(csr_wrdata[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_18),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[18] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[18] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[19] (
	.clk(clk),
	.d(csr_wrdata[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_19),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[19] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[19] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[19] (
	.clk(clk),
	.d(csr_wrdata[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_19),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[19] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[19] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[19] (
	.clk(clk),
	.d(csr_wrdata[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_19),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[19] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[19] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[20] (
	.clk(clk),
	.d(csr_wrdata[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_20),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[20] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[20] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[20] (
	.clk(clk),
	.d(csr_wrdata[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_20),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[20] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[20] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[20] (
	.clk(clk),
	.d(csr_wrdata[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_20),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[20] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[20] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[21] (
	.clk(clk),
	.d(csr_wrdata[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_21),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[21] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[21] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[21] (
	.clk(clk),
	.d(csr_wrdata[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_21),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[21] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[21] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[21] (
	.clk(clk),
	.d(csr_wrdata[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_21),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[21] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[21] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[22] (
	.clk(clk),
	.d(csr_wrdata[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_22),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[22] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[22] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[22] (
	.clk(clk),
	.d(csr_wrdata[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_22),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[22] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[22] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[22] (
	.clk(clk),
	.d(csr_wrdata[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_22),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[22] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[22] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[23] (
	.clk(clk),
	.d(csr_wrdata[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_23),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[23] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[23] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[23] (
	.clk(clk),
	.d(csr_wrdata[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_23),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[23] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[23] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[23] (
	.clk(clk),
	.d(csr_wrdata[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_23),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[23] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[23] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[24] (
	.clk(clk),
	.d(csr_wrdata[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_24),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[24] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[24] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[24] (
	.clk(clk),
	.d(csr_wrdata[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_24),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[24] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[24] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[24] (
	.clk(clk),
	.d(csr_wrdata[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_24),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[24] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[24] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[25] (
	.clk(clk),
	.d(csr_wrdata[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_25),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[25] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[25] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[25] (
	.clk(clk),
	.d(csr_wrdata[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_25),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[25] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[25] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[25] (
	.clk(clk),
	.d(csr_wrdata[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_25),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[25] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[25] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[26] (
	.clk(clk),
	.d(csr_wrdata[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_26),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[26] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[26] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[26] (
	.clk(clk),
	.d(csr_wrdata[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_26),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[26] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[26] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[26] (
	.clk(clk),
	.d(csr_wrdata[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_26),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[26] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[26] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[27] (
	.clk(clk),
	.d(csr_wrdata[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_27),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[27] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[27] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[27] (
	.clk(clk),
	.d(csr_wrdata[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_27),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[27] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[27] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[27] (
	.clk(clk),
	.d(csr_wrdata[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_27),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[27] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[27] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[28] (
	.clk(clk),
	.d(csr_wrdata[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_28),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[28] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[28] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[28] (
	.clk(clk),
	.d(csr_wrdata[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_28),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[28] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[28] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[28] (
	.clk(clk),
	.d(csr_wrdata[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_28),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[28] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[28] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[29] (
	.clk(clk),
	.d(csr_wrdata[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_29),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[29] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[29] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[29] (
	.clk(clk),
	.d(csr_wrdata[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_29),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[29] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[29] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[29] (
	.clk(clk),
	.d(csr_wrdata[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_29),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[29] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[29] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[30] (
	.clk(clk),
	.d(csr_wrdata[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_30),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[30] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[30] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[30] (
	.clk(clk),
	.d(csr_wrdata[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_30),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[30] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[30] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[30] (
	.clk(clk),
	.d(csr_wrdata[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_30),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[30] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[30] .power_up = "low";

dffeas \csr_flash_cmd_addr_data[31] (
	.clk(clk),
	.d(csr_wrdata[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_addr~combout ),
	.q(csr_flash_cmd_addr_data_31),
	.prn(vcc));
defparam \csr_flash_cmd_addr_data[31] .is_wysiwyg = "true";
defparam \csr_flash_cmd_addr_data[31] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_0_data[31] (
	.clk(clk),
	.d(csr_wrdata[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_0~combout ),
	.q(csr_flash_cmd_wr_data_0_data_31),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_0_data[31] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_0_data[31] .power_up = "low";

dffeas \csr_flash_cmd_wr_data_1_data[31] (
	.clk(clk),
	.d(csr_wrdata[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_wr_data_1~combout ),
	.q(csr_flash_cmd_wr_data_1_data_31),
	.prn(vcc));
defparam \csr_flash_cmd_wr_data_1_data[31] .is_wysiwyg = "true";
defparam \csr_flash_cmd_wr_data_1_data[31] .power_up = "low";

dffeas \state.ST_WAIT_RSP (
	.clk(clk),
	.d(\Selector36~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stateST_WAIT_RSP),
	.prn(vcc));
defparam \state.ST_WAIT_RSP .is_wysiwyg = "true";
defparam \state.ST_WAIT_RSP .power_up = "low";

dffeas \state.ST_SEND_HEADER (
	.clk(clk),
	.d(\Selector33~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stateST_SEND_HEADER),
	.prn(vcc));
defparam \state.ST_SEND_HEADER .is_wysiwyg = "true";
defparam \state.ST_SEND_HEADER .power_up = "low";

dffeas \state.ST_SEND_DATA_1 (
	.clk(clk),
	.d(\Selector35~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sink1_ready),
	.q(stateST_SEND_DATA_1),
	.prn(vcc));
defparam \state.ST_SEND_DATA_1 .is_wysiwyg = "true";
defparam \state.ST_SEND_DATA_1 .power_up = "low";

dffeas \state.ST_SEND_DATA_0 (
	.clk(clk),
	.d(Selector34),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sink1_ready),
	.q(stateST_SEND_DATA_0),
	.prn(vcc));
defparam \state.ST_SEND_DATA_0 .is_wysiwyg = "true";
defparam \state.ST_SEND_DATA_0 .power_up = "low";

dffeas has_data_in(
	.clk(clk),
	.d(\has_data_in~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(has_data_in1),
	.prn(vcc));
defparam has_data_in.is_wysiwyg = "true";
defparam has_data_in.power_up = "low";

dffeas more_than_4bytes_data(
	.clk(clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(more_than_4bytes_data1),
	.prn(vcc));
defparam more_than_4bytes_data.is_wysiwyg = "true";
defparam more_than_4bytes_data.power_up = "low";

cycloneive_lcell_comb \Selector34~0 (
	.dataa(stateST_SEND_HEADER),
	.datab(has_data_in1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(Selector34),
	.cout());
defparam \Selector34~0 .lut_mask = 16'h8888;
defparam \Selector34~0 .sum_lutc_input = "datac";

dffeas has_data_out(
	.clk(clk),
	.d(\has_data_out~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(has_data_out1),
	.prn(vcc));
defparam has_data_out.is_wysiwyg = "true";
defparam has_data_out.power_up = "low";

dffeas \numb_data[0] (
	.clk(clk),
	.d(\numb_data[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(numb_data_0),
	.prn(vcc));
defparam \numb_data[0] .is_wysiwyg = "true";
defparam \numb_data[0] .power_up = "low";

dffeas \numb_data[1] (
	.clk(clk),
	.d(\csr_flash_cmd_setting_data[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(numb_data_1),
	.prn(vcc));
defparam \numb_data[1] .is_wysiwyg = "true";
defparam \numb_data[1] .power_up = "low";

dffeas \numb_data[3] (
	.clk(clk),
	.d(\csr_flash_cmd_setting_data[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(numb_data_3),
	.prn(vcc));
defparam \numb_data[3] .is_wysiwyg = "true";
defparam \numb_data[3] .power_up = "low";

dffeas \numb_data[2] (
	.clk(clk),
	.d(\csr_flash_cmd_setting_data[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(numb_data_2),
	.prn(vcc));
defparam \numb_data[2] .is_wysiwyg = "true";
defparam \numb_data[2] .power_up = "low";

dffeas has_addr(
	.clk(clk),
	.d(\Equal13~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(has_addr1),
	.prn(vcc));
defparam has_addr.is_wysiwyg = "true";
defparam has_addr.power_up = "low";

dffeas \numb_dummy[0] (
	.clk(clk),
	.d(\csr_flash_cmd_setting_data[16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(numb_dummy_0),
	.prn(vcc));
defparam \numb_dummy[0] .is_wysiwyg = "true";
defparam \numb_dummy[0] .power_up = "low";

dffeas \numb_dummy[4] (
	.clk(clk),
	.d(\csr_flash_cmd_setting_data[20]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(numb_dummy_4),
	.prn(vcc));
defparam \numb_dummy[4] .is_wysiwyg = "true";
defparam \numb_dummy[4] .power_up = "low";

dffeas \numb_dummy[3] (
	.clk(clk),
	.d(\csr_flash_cmd_setting_data[19]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(numb_dummy_3),
	.prn(vcc));
defparam \numb_dummy[3] .is_wysiwyg = "true";
defparam \numb_dummy[3] .power_up = "low";

dffeas \numb_dummy[2] (
	.clk(clk),
	.d(\csr_flash_cmd_setting_data[18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(numb_dummy_2),
	.prn(vcc));
defparam \numb_dummy[2] .is_wysiwyg = "true";
defparam \numb_dummy[2] .power_up = "low";

dffeas \numb_dummy[1] (
	.clk(clk),
	.d(\csr_flash_cmd_setting_data[17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(numb_dummy_1),
	.prn(vcc));
defparam \numb_dummy[1] .is_wysiwyg = "true";
defparam \numb_dummy[1] .power_up = "low";

dffeas is_4bytes_addr(
	.clk(clk),
	.d(\Equal14~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(is_4bytes_addr1),
	.prn(vcc));
defparam is_4bytes_addr.is_wysiwyg = "true";
defparam is_4bytes_addr.power_up = "low";

dffeas \opcode[0] (
	.clk(clk),
	.d(\opcode[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(opcode_0),
	.prn(vcc));
defparam \opcode[0] .is_wysiwyg = "true";
defparam \opcode[0] .power_up = "low";

dffeas \opcode[4] (
	.clk(clk),
	.d(\csr_flash_cmd_setting_data[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(opcode_4),
	.prn(vcc));
defparam \opcode[4] .is_wysiwyg = "true";
defparam \opcode[4] .power_up = "low";

dffeas \opcode[2] (
	.clk(clk),
	.d(\opcode[2]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(opcode_2),
	.prn(vcc));
defparam \opcode[2] .is_wysiwyg = "true";
defparam \opcode[2] .power_up = "low";

dffeas \opcode[1] (
	.clk(clk),
	.d(\csr_flash_cmd_setting_data[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(opcode_1),
	.prn(vcc));
defparam \opcode[1] .is_wysiwyg = "true";
defparam \opcode[1] .power_up = "low";

dffeas \opcode[3] (
	.clk(clk),
	.d(\csr_flash_cmd_setting_data[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(opcode_3),
	.prn(vcc));
defparam \opcode[3] .is_wysiwyg = "true";
defparam \opcode[3] .power_up = "low";

dffeas \opcode[5] (
	.clk(clk),
	.d(\csr_flash_cmd_setting_data[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(opcode_5),
	.prn(vcc));
defparam \opcode[5] .is_wysiwyg = "true";
defparam \opcode[5] .power_up = "low";

dffeas \opcode[6] (
	.clk(clk),
	.d(\csr_flash_cmd_setting_data[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(opcode_6),
	.prn(vcc));
defparam \opcode[6] .is_wysiwyg = "true";
defparam \opcode[6] .power_up = "low";

dffeas \opcode[7] (
	.clk(clk),
	.d(\csr_flash_cmd_setting_data[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(opcode_7),
	.prn(vcc));
defparam \opcode[7] .is_wysiwyg = "true";
defparam \opcode[7] .power_up = "low";

dffeas has_dummy(
	.clk(clk),
	.d(\Equal15~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(has_dummy1),
	.prn(vcc));
defparam has_dummy.is_wysiwyg = "true";
defparam has_dummy.power_up = "low";

cycloneive_lcell_comb \rdata_comb[0]~2 (
	.dataa(avl_csr_address_1),
	.datab(csr_rd_inst_data_0),
	.datac(avl_csr_address_0),
	.datad(csr_op_protocol_data_0),
	.cin(gnd),
	.combout(\rdata_comb[0]~2_combout ),
	.cout());
defparam \rdata_comb[0]~2 .lut_mask = 16'hB5B0;
defparam \rdata_comb[0]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \csr_flash_cmd_setting_data[0]~0 (
	.dataa(csr_wrdata[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\csr_flash_cmd_setting_data[0]~0_combout ),
	.cout());
defparam \csr_flash_cmd_setting_data[0]~0 .lut_mask = 16'h5555;
defparam \csr_flash_cmd_setting_data[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_csr_control~0 (
	.dataa(avl_csr_write),
	.datab(csr_waitrequest1),
	.datac(avl_csr_address_4),
	.datad(avl_csr_address_5),
	.cin(gnd),
	.combout(\wr_csr_control~0_combout ),
	.cout());
defparam \wr_csr_control~0 .lut_mask = 16'h0002;
defparam \wr_csr_control~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_csr_op_protocol~0 (
	.dataa(avl_csr_address_2),
	.datab(\wr_csr_control~0_combout ),
	.datac(gnd),
	.datad(avl_csr_address_3),
	.cin(gnd),
	.combout(\wr_csr_op_protocol~0_combout ),
	.cout());
defparam \wr_csr_op_protocol~0 .lut_mask = 16'h0088;
defparam \wr_csr_op_protocol~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb wr_csr_flash_cmd_setting(
	.dataa(avl_csr_address_1),
	.datab(avl_csr_address_0),
	.datac(\wr_csr_op_protocol~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_csr_flash_cmd_setting~combout ),
	.cout());
defparam wr_csr_flash_cmd_setting.lut_mask = 16'h8080;
defparam wr_csr_flash_cmd_setting.sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[0] (
	.clk(clk),
	.d(\csr_flash_cmd_setting_data[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[0]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[0] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[0] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[0]~3 (
	.dataa(csr_wr_inst_data_0),
	.datab(avl_csr_address_1),
	.datac(\rdata_comb[0]~2_combout ),
	.datad(\csr_flash_cmd_setting_data[0]~q ),
	.cin(gnd),
	.combout(\rdata_comb[0]~3_combout ),
	.cout());
defparam \rdata_comb[0]~3 .lut_mask = 16'h38F8;
defparam \rdata_comb[0]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \avl_rddata_local[3]~2 (
	.dataa(avl_csr_address_2),
	.datab(avl_csr_address_0),
	.datac(avl_csr_address_1),
	.datad(avl_csr_address_3),
	.cin(gnd),
	.combout(\avl_rddata_local[3]~2_combout ),
	.cout());
defparam \avl_rddata_local[3]~2 .lut_mask = 16'h08AA;
defparam \avl_rddata_local[3]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \avl_rddata_local[3]~3 (
	.dataa(avl_csr_address_1),
	.datab(gnd),
	.datac(gnd),
	.datad(avl_csr_address_2),
	.cin(gnd),
	.combout(\avl_rddata_local[3]~3_combout ),
	.cout());
defparam \avl_rddata_local[3]~3 .lut_mask = 16'h00AA;
defparam \avl_rddata_local[3]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_data_cnt~1 (
	.dataa(\read_data_cnt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(stateST_IDLE),
	.cin(gnd),
	.combout(\read_data_cnt~1_combout ),
	.cout());
defparam \read_data_cnt~1 .lut_mask = 16'h5500;
defparam \read_data_cnt~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \read_data_cnt[0]~2 (
	.dataa(sink_ready),
	.datab(out_valid),
	.datac(stateST_SEND_DUMMY_RSP),
	.datad(stateST_IDLE),
	.cin(gnd),
	.combout(\read_data_cnt[0]~2_combout ),
	.cout());
defparam \read_data_cnt[0]~2 .lut_mask = 16'hA8FF;
defparam \read_data_cnt[0]~2 .sum_lutc_input = "datac";

dffeas \read_data_cnt[0] (
	.clk(clk),
	.d(\read_data_cnt~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_cnt[0]~2_combout ),
	.q(\read_data_cnt[0]~q ),
	.prn(vcc));
defparam \read_data_cnt[0] .is_wysiwyg = "true";
defparam \read_data_cnt[0] .power_up = "low";

cycloneive_lcell_comb \read_data_cnt~3 (
	.dataa(stateST_IDLE),
	.datab(gnd),
	.datac(\read_data_cnt[0]~q ),
	.datad(\read_data_cnt[1]~q ),
	.cin(gnd),
	.combout(\read_data_cnt~3_combout ),
	.cout());
defparam \read_data_cnt~3 .lut_mask = 16'h0AA0;
defparam \read_data_cnt~3 .sum_lutc_input = "datac";

dffeas \read_data_cnt[1] (
	.clk(clk),
	.d(\read_data_cnt~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_cnt[0]~2_combout ),
	.q(\read_data_cnt[1]~q ),
	.prn(vcc));
defparam \read_data_cnt[1] .is_wysiwyg = "true";
defparam \read_data_cnt[1] .power_up = "low";

cycloneive_lcell_comb \csr_flash_cmd_rd_data_0_data[0]~0 (
	.dataa(stateST_WAIT_RSP),
	.datab(gnd),
	.datac(\read_data_cnt[0]~q ),
	.datad(\read_data_cnt[1]~q ),
	.cin(gnd),
	.combout(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.cout());
defparam \csr_flash_cmd_rd_data_0_data[0]~0 .lut_mask = 16'h000A;
defparam \csr_flash_cmd_rd_data_0_data[0]~0 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_0_data[0] (
	.clk(clk),
	.d(out_rsp_data_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[0]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[0] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[0] .power_up = "low";

cycloneive_lcell_comb \avl_rddata_local[3]~4 (
	.dataa(avl_csr_address_2),
	.datab(avl_csr_address_1),
	.datac(avl_csr_address_0),
	.datad(gnd),
	.cin(gnd),
	.combout(\avl_rddata_local[3]~4_combout ),
	.cout());
defparam \avl_rddata_local[3]~4 .lut_mask = 16'hEAEA;
defparam \avl_rddata_local[3]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[0]~4 (
	.dataa(\avl_rddata_local[3]~3_combout ),
	.datab(\csr_flash_cmd_rd_data_0_data[0]~q ),
	.datac(\avl_rddata_local[3]~4_combout ),
	.datad(csr_flash_cmd_addr_data_0),
	.cin(gnd),
	.combout(\rdata_comb[0]~4_combout ),
	.cout());
defparam \rdata_comb[0]~4 .lut_mask = 16'hE5E0;
defparam \rdata_comb[0]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[0]~5 (
	.dataa(csr_flash_cmd_wr_data_0_data_0),
	.datab(\avl_rddata_local[3]~3_combout ),
	.datac(\rdata_comb[0]~4_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_0),
	.cin(gnd),
	.combout(\rdata_comb[0]~5_combout ),
	.cout());
defparam \rdata_comb[0]~5 .lut_mask = 16'hF838;
defparam \rdata_comb[0]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[0]~6 (
	.dataa(avl_csr_address_1),
	.datab(csr_clk_baud_rate_data_0),
	.datac(avl_csr_address_0),
	.datad(csr_control_data_0),
	.cin(gnd),
	.combout(\rdata_comb[0]~6_combout ),
	.cout());
defparam \rdata_comb[0]~6 .lut_mask = 16'hE0E5;
defparam \rdata_comb[0]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[0]~7 (
	.dataa(csr_delay_setting_data_0),
	.datab(avl_csr_address_1),
	.datac(\rdata_comb[0]~6_combout ),
	.datad(csr_rd_capturing_data_0),
	.cin(gnd),
	.combout(\rdata_comb[0]~7_combout ),
	.cout());
defparam \rdata_comb[0]~7 .lut_mask = 16'hF838;
defparam \rdata_comb[0]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[0]~8 (
	.dataa(\avl_rddata_local[3]~2_combout ),
	.datab(\rdata_comb[0]~5_combout ),
	.datac(avl_csr_address_3),
	.datad(\rdata_comb[0]~7_combout ),
	.cin(gnd),
	.combout(\rdata_comb[0]~8_combout ),
	.cout());
defparam \rdata_comb[0]~8 .lut_mask = 16'hE5E0;
defparam \rdata_comb[0]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \csr_flash_cmd_rd_data_1_data[0]~0 (
	.dataa(stateST_WAIT_RSP),
	.datab(\read_data_cnt[0]~q ),
	.datac(gnd),
	.datad(\read_data_cnt[1]~q ),
	.cin(gnd),
	.combout(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.cout());
defparam \csr_flash_cmd_rd_data_1_data[0]~0 .lut_mask = 16'h0088;
defparam \csr_flash_cmd_rd_data_1_data[0]~0 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[0] (
	.clk(clk),
	.d(out_rsp_data_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[0]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[0] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[0] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[0]~9 (
	.dataa(\rdata_comb[0]~3_combout ),
	.datab(\avl_rddata_local[3]~2_combout ),
	.datac(\rdata_comb[0]~8_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[0]~q ),
	.cin(gnd),
	.combout(\rdata_comb[0]~9_combout ),
	.cout());
defparam \rdata_comb[0]~9 .lut_mask = 16'hF838;
defparam \rdata_comb[0]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[4]~10 (
	.dataa(avl_csr_read),
	.datab(gnd),
	.datac(avl_csr_address_4),
	.datad(avl_csr_address_5),
	.cin(gnd),
	.combout(\rdata_comb[4]~10_combout ),
	.cout());
defparam \rdata_comb[4]~10 .lut_mask = 16'h000A;
defparam \rdata_comb[4]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \avl_rddata_local[3]~5 (
	.dataa(avl_csr_address_3),
	.datab(avl_csr_address_1),
	.datac(avl_csr_address_2),
	.datad(avl_csr_address_0),
	.cin(gnd),
	.combout(\avl_rddata_local[3]~5_combout ),
	.cout());
defparam \avl_rddata_local[3]~5 .lut_mask = 16'h8082;
defparam \avl_rddata_local[3]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[0]~11 (
	.dataa(\rdata_comb[0]~9_combout ),
	.datab(\rdata_comb[4]~10_combout ),
	.datac(gnd),
	.datad(\avl_rddata_local[3]~5_combout ),
	.cin(gnd),
	.combout(\rdata_comb[0]~11_combout ),
	.cout());
defparam \rdata_comb[0]~11 .lut_mask = 16'h0088;
defparam \rdata_comb[0]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[1]~12 (
	.dataa(avl_csr_address_1),
	.datab(csr_rd_inst_data_1),
	.datac(avl_csr_address_0),
	.datad(csr_op_protocol_data_1),
	.cin(gnd),
	.combout(\rdata_comb[1]~12_combout ),
	.cout());
defparam \rdata_comb[1]~12 .lut_mask = 16'hB5B0;
defparam \rdata_comb[1]~12 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[1] (
	.clk(clk),
	.d(csr_wrdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[1]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[1] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[1] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[1]~13 (
	.dataa(csr_wr_inst_data_1),
	.datab(avl_csr_address_1),
	.datac(\rdata_comb[1]~12_combout ),
	.datad(\csr_flash_cmd_setting_data[1]~q ),
	.cin(gnd),
	.combout(\rdata_comb[1]~13_combout ),
	.cout());
defparam \rdata_comb[1]~13 .lut_mask = 16'hF434;
defparam \rdata_comb[1]~13 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_0_data[1] (
	.clk(clk),
	.d(out_rsp_data_1),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[1]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[1] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[1] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[1]~14 (
	.dataa(\avl_rddata_local[3]~4_combout ),
	.datab(csr_flash_cmd_wr_data_0_data_1),
	.datac(\avl_rddata_local[3]~3_combout ),
	.datad(csr_flash_cmd_addr_data_1),
	.cin(gnd),
	.combout(\rdata_comb[1]~14_combout ),
	.cout());
defparam \rdata_comb[1]~14 .lut_mask = 16'hE5E0;
defparam \rdata_comb[1]~14 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[1]~15 (
	.dataa(\csr_flash_cmd_rd_data_0_data[1]~q ),
	.datab(\avl_rddata_local[3]~4_combout ),
	.datac(\rdata_comb[1]~14_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_1),
	.cin(gnd),
	.combout(\rdata_comb[1]~15_combout ),
	.cout());
defparam \rdata_comb[1]~15 .lut_mask = 16'hF838;
defparam \rdata_comb[1]~15 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_csr_control~1 (
	.dataa(\wr_csr_control~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(avl_csr_address_2),
	.cin(gnd),
	.combout(\wr_csr_control~1_combout ),
	.cout());
defparam \wr_csr_control~1 .lut_mask = 16'h00AA;
defparam \wr_csr_control~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb wr_csr_control(
	.dataa(\wr_csr_control~1_combout ),
	.datab(avl_csr_address_1),
	.datac(avl_csr_address_0),
	.datad(avl_csr_address_3),
	.cin(gnd),
	.combout(\wr_csr_control~combout ),
	.cout());
defparam wr_csr_control.lut_mask = 16'h0002;
defparam wr_csr_control.sum_lutc_input = "datac";

dffeas \csr_control_data[1] (
	.clk(clk),
	.d(csr_wrdata[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[1]~q ),
	.prn(vcc));
defparam \csr_control_data[1] .is_wysiwyg = "true";
defparam \csr_control_data[1] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[1]~16 (
	.dataa(avl_csr_address_1),
	.datab(csr_clk_baud_rate_data_1),
	.datac(avl_csr_address_0),
	.datad(\csr_control_data[1]~q ),
	.cin(gnd),
	.combout(\rdata_comb[1]~16_combout ),
	.cout());
defparam \rdata_comb[1]~16 .lut_mask = 16'hE5E0;
defparam \rdata_comb[1]~16 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[1]~17 (
	.dataa(csr_delay_setting_data_1),
	.datab(avl_csr_address_1),
	.datac(\rdata_comb[1]~16_combout ),
	.datad(csr_rd_capturing_data_1),
	.cin(gnd),
	.combout(\rdata_comb[1]~17_combout ),
	.cout());
defparam \rdata_comb[1]~17 .lut_mask = 16'hF838;
defparam \rdata_comb[1]~17 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[1]~18 (
	.dataa(\avl_rddata_local[3]~2_combout ),
	.datab(\rdata_comb[1]~15_combout ),
	.datac(avl_csr_address_3),
	.datad(\rdata_comb[1]~17_combout ),
	.cin(gnd),
	.combout(\rdata_comb[1]~18_combout ),
	.cout());
defparam \rdata_comb[1]~18 .lut_mask = 16'hE5E0;
defparam \rdata_comb[1]~18 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[1] (
	.clk(clk),
	.d(out_rsp_data_1),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[1]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[1] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[1] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[1]~19 (
	.dataa(\rdata_comb[1]~13_combout ),
	.datab(\avl_rddata_local[3]~2_combout ),
	.datac(\rdata_comb[1]~18_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[1]~q ),
	.cin(gnd),
	.combout(\rdata_comb[1]~19_combout ),
	.cout());
defparam \rdata_comb[1]~19 .lut_mask = 16'hF838;
defparam \rdata_comb[1]~19 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[1]~20 (
	.dataa(\rdata_comb[4]~10_combout ),
	.datab(\rdata_comb[1]~19_combout ),
	.datac(gnd),
	.datad(\avl_rddata_local[3]~5_combout ),
	.cin(gnd),
	.combout(\rdata_comb[1]~20_combout ),
	.cout());
defparam \rdata_comb[1]~20 .lut_mask = 16'h0088;
defparam \rdata_comb[1]~20 .sum_lutc_input = "datac";

cycloneive_lcell_comb wr_csr_op_protocol(
	.dataa(\wr_csr_op_protocol~0_combout ),
	.datab(gnd),
	.datac(avl_csr_address_1),
	.datad(avl_csr_address_0),
	.cin(gnd),
	.combout(\wr_csr_op_protocol~combout ),
	.cout());
defparam wr_csr_op_protocol.lut_mask = 16'h000A;
defparam wr_csr_op_protocol.sum_lutc_input = "datac";

dffeas \csr_op_protocol_data[2] (
	.clk(clk),
	.d(csr_wrdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(\csr_op_protocol_data[2]~q ),
	.prn(vcc));
defparam \csr_op_protocol_data[2] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[2] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[2]~21 (
	.dataa(avl_csr_address_1),
	.datab(csr_rd_inst_data_2),
	.datac(avl_csr_address_0),
	.datad(\csr_op_protocol_data[2]~q ),
	.cin(gnd),
	.combout(\rdata_comb[2]~21_combout ),
	.cout());
defparam \rdata_comb[2]~21 .lut_mask = 16'hE5E0;
defparam \rdata_comb[2]~21 .sum_lutc_input = "datac";

cycloneive_lcell_comb \csr_flash_cmd_setting_data[2]~1 (
	.dataa(csr_wrdata[2]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\csr_flash_cmd_setting_data[2]~1_combout ),
	.cout());
defparam \csr_flash_cmd_setting_data[2]~1 .lut_mask = 16'h5555;
defparam \csr_flash_cmd_setting_data[2]~1 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[2] (
	.clk(clk),
	.d(\csr_flash_cmd_setting_data[2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[2]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[2] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[2] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[2]~22 (
	.dataa(csr_wr_inst_data_2),
	.datab(avl_csr_address_1),
	.datac(\rdata_comb[2]~21_combout ),
	.datad(\csr_flash_cmd_setting_data[2]~q ),
	.cin(gnd),
	.combout(\rdata_comb[2]~22_combout ),
	.cout());
defparam \rdata_comb[2]~22 .lut_mask = 16'h38F8;
defparam \rdata_comb[2]~22 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_0_data[2] (
	.clk(clk),
	.d(out_rsp_data_2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[2]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[2] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[2] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[2]~23 (
	.dataa(\avl_rddata_local[3]~3_combout ),
	.datab(\csr_flash_cmd_rd_data_0_data[2]~q ),
	.datac(\avl_rddata_local[3]~4_combout ),
	.datad(csr_flash_cmd_addr_data_2),
	.cin(gnd),
	.combout(\rdata_comb[2]~23_combout ),
	.cout());
defparam \rdata_comb[2]~23 .lut_mask = 16'hE5E0;
defparam \rdata_comb[2]~23 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[2]~24 (
	.dataa(csr_flash_cmd_wr_data_0_data_2),
	.datab(\avl_rddata_local[3]~3_combout ),
	.datac(\rdata_comb[2]~23_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_2),
	.cin(gnd),
	.combout(\rdata_comb[2]~24_combout ),
	.cout());
defparam \rdata_comb[2]~24 .lut_mask = 16'hF838;
defparam \rdata_comb[2]~24 .sum_lutc_input = "datac";

dffeas \csr_control_data[2] (
	.clk(clk),
	.d(csr_wrdata[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[2]~q ),
	.prn(vcc));
defparam \csr_control_data[2] .is_wysiwyg = "true";
defparam \csr_control_data[2] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[2]~25 (
	.dataa(avl_csr_address_1),
	.datab(csr_clk_baud_rate_data_2),
	.datac(avl_csr_address_0),
	.datad(\csr_control_data[2]~q ),
	.cin(gnd),
	.combout(\rdata_comb[2]~25_combout ),
	.cout());
defparam \rdata_comb[2]~25 .lut_mask = 16'hE5E0;
defparam \rdata_comb[2]~25 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[2]~26 (
	.dataa(csr_delay_setting_data_2),
	.datab(avl_csr_address_1),
	.datac(\rdata_comb[2]~25_combout ),
	.datad(csr_rd_capturing_data_2),
	.cin(gnd),
	.combout(\rdata_comb[2]~26_combout ),
	.cout());
defparam \rdata_comb[2]~26 .lut_mask = 16'hF838;
defparam \rdata_comb[2]~26 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[2]~27 (
	.dataa(\avl_rddata_local[3]~2_combout ),
	.datab(\rdata_comb[2]~24_combout ),
	.datac(avl_csr_address_3),
	.datad(\rdata_comb[2]~26_combout ),
	.cin(gnd),
	.combout(\rdata_comb[2]~27_combout ),
	.cout());
defparam \rdata_comb[2]~27 .lut_mask = 16'hE5E0;
defparam \rdata_comb[2]~27 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[2] (
	.clk(clk),
	.d(out_rsp_data_2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[2]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[2] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[2] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[2]~28 (
	.dataa(\rdata_comb[2]~22_combout ),
	.datab(\avl_rddata_local[3]~2_combout ),
	.datac(\rdata_comb[2]~27_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[2]~q ),
	.cin(gnd),
	.combout(\rdata_comb[2]~28_combout ),
	.cout());
defparam \rdata_comb[2]~28 .lut_mask = 16'hF838;
defparam \rdata_comb[2]~28 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[2]~29 (
	.dataa(\rdata_comb[4]~10_combout ),
	.datab(\rdata_comb[2]~28_combout ),
	.datac(gnd),
	.datad(\avl_rddata_local[3]~5_combout ),
	.cin(gnd),
	.combout(\rdata_comb[2]~29_combout ),
	.cout());
defparam \rdata_comb[2]~29 .lut_mask = 16'h0088;
defparam \rdata_comb[2]~29 .sum_lutc_input = "datac";

dffeas \csr_op_protocol_data[3] (
	.clk(clk),
	.d(csr_wrdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(\csr_op_protocol_data[3]~q ),
	.prn(vcc));
defparam \csr_op_protocol_data[3] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[3] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[3]~30 (
	.dataa(avl_csr_address_1),
	.datab(csr_rd_inst_data_3),
	.datac(avl_csr_address_0),
	.datad(\csr_op_protocol_data[3]~q ),
	.cin(gnd),
	.combout(\rdata_comb[3]~30_combout ),
	.cout());
defparam \rdata_comb[3]~30 .lut_mask = 16'hE5E0;
defparam \rdata_comb[3]~30 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[3] (
	.clk(clk),
	.d(csr_wrdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[3]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[3] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[3] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[3]~31 (
	.dataa(csr_wr_inst_data_3),
	.datab(avl_csr_address_1),
	.datac(\rdata_comb[3]~30_combout ),
	.datad(\csr_flash_cmd_setting_data[3]~q ),
	.cin(gnd),
	.combout(\rdata_comb[3]~31_combout ),
	.cout());
defparam \rdata_comb[3]~31 .lut_mask = 16'hF838;
defparam \rdata_comb[3]~31 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_0_data[3] (
	.clk(clk),
	.d(out_rsp_data_3),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[3]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[3] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[3] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[3]~32 (
	.dataa(\avl_rddata_local[3]~4_combout ),
	.datab(csr_flash_cmd_wr_data_0_data_3),
	.datac(\avl_rddata_local[3]~3_combout ),
	.datad(csr_flash_cmd_addr_data_3),
	.cin(gnd),
	.combout(\rdata_comb[3]~32_combout ),
	.cout());
defparam \rdata_comb[3]~32 .lut_mask = 16'hE5E0;
defparam \rdata_comb[3]~32 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[3]~33 (
	.dataa(\csr_flash_cmd_rd_data_0_data[3]~q ),
	.datab(\avl_rddata_local[3]~4_combout ),
	.datac(\rdata_comb[3]~32_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_3),
	.cin(gnd),
	.combout(\rdata_comb[3]~33_combout ),
	.cout());
defparam \rdata_comb[3]~33 .lut_mask = 16'hF838;
defparam \rdata_comb[3]~33 .sum_lutc_input = "datac";

dffeas \csr_control_data[3] (
	.clk(clk),
	.d(csr_wrdata[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[3]~q ),
	.prn(vcc));
defparam \csr_control_data[3] .is_wysiwyg = "true";
defparam \csr_control_data[3] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[3]~34 (
	.dataa(avl_csr_address_1),
	.datab(csr_clk_baud_rate_data_3),
	.datac(avl_csr_address_0),
	.datad(\csr_control_data[3]~q ),
	.cin(gnd),
	.combout(\rdata_comb[3]~34_combout ),
	.cout());
defparam \rdata_comb[3]~34 .lut_mask = 16'hE5E0;
defparam \rdata_comb[3]~34 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[3]~35 (
	.dataa(csr_delay_setting_data_3),
	.datab(avl_csr_address_1),
	.datac(\rdata_comb[3]~34_combout ),
	.datad(csr_rd_capturing_data_3),
	.cin(gnd),
	.combout(\rdata_comb[3]~35_combout ),
	.cout());
defparam \rdata_comb[3]~35 .lut_mask = 16'hF838;
defparam \rdata_comb[3]~35 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[3]~36 (
	.dataa(\avl_rddata_local[3]~2_combout ),
	.datab(\rdata_comb[3]~33_combout ),
	.datac(avl_csr_address_3),
	.datad(\rdata_comb[3]~35_combout ),
	.cin(gnd),
	.combout(\rdata_comb[3]~36_combout ),
	.cout());
defparam \rdata_comb[3]~36 .lut_mask = 16'hE5E0;
defparam \rdata_comb[3]~36 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[3] (
	.clk(clk),
	.d(out_rsp_data_3),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[3]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[3] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[3] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[3]~37 (
	.dataa(\rdata_comb[3]~31_combout ),
	.datab(\avl_rddata_local[3]~2_combout ),
	.datac(\rdata_comb[3]~36_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[3]~q ),
	.cin(gnd),
	.combout(\rdata_comb[3]~37_combout ),
	.cout());
defparam \rdata_comb[3]~37 .lut_mask = 16'hF838;
defparam \rdata_comb[3]~37 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[3]~38 (
	.dataa(\rdata_comb[4]~10_combout ),
	.datab(\rdata_comb[3]~37_combout ),
	.datac(gnd),
	.datad(\avl_rddata_local[3]~5_combout ),
	.cin(gnd),
	.combout(\rdata_comb[3]~38_combout ),
	.cout());
defparam \rdata_comb[3]~38 .lut_mask = 16'h0088;
defparam \rdata_comb[3]~38 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector27~0 (
	.dataa(csr_wr_inst_data_4),
	.datab(csr_delay_setting_data_4),
	.datac(avl_csr_address_2),
	.datad(avl_csr_address_0),
	.cin(gnd),
	.combout(\Selector27~0_combout ),
	.cout());
defparam \Selector27~0 .lut_mask = 16'h00AC;
defparam \Selector27~0 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[4] (
	.clk(clk),
	.d(csr_wrdata[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[4]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[4] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[4] .power_up = "low";

cycloneive_lcell_comb \Selector27~1 (
	.dataa(\Selector27~0_combout ),
	.datab(avl_csr_address_0),
	.datac(avl_csr_address_2),
	.datad(\csr_flash_cmd_setting_data[4]~q ),
	.cin(gnd),
	.combout(\Selector27~1_combout ),
	.cout());
defparam \Selector27~1 .lut_mask = 16'hEAAA;
defparam \Selector27~1 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[4] (
	.clk(clk),
	.d(out_rsp_data_4),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[4]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[4] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[4] .power_up = "low";

dffeas \csr_flash_cmd_rd_data_0_data[4] (
	.clk(clk),
	.d(out_rsp_data_4),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[4]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[4] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[4] .power_up = "low";

cycloneive_lcell_comb \Selector27~2 (
	.dataa(avl_csr_address_2),
	.datab(\csr_flash_cmd_rd_data_1_data[4]~q ),
	.datac(\csr_flash_cmd_rd_data_0_data[4]~q ),
	.datad(avl_csr_address_0),
	.cin(gnd),
	.combout(\Selector27~2_combout ),
	.cout());
defparam \Selector27~2 .lut_mask = 16'h88A0;
defparam \Selector27~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector27~3 (
	.dataa(\Selector27~2_combout ),
	.datab(avl_csr_address_0),
	.datac(csr_flash_cmd_addr_data_4),
	.datad(avl_csr_address_2),
	.cin(gnd),
	.combout(\Selector27~3_combout ),
	.cout());
defparam \Selector27~3 .lut_mask = 16'hAAEA;
defparam \Selector27~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector27~4 (
	.dataa(avl_csr_address_2),
	.datab(csr_clk_baud_rate_data_4),
	.datac(avl_csr_address_0),
	.datad(csr_control_data_4),
	.cin(gnd),
	.combout(\Selector27~4_combout ),
	.cout());
defparam \Selector27~4 .lut_mask = 16'hB5B0;
defparam \Selector27~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector27~5 (
	.dataa(csr_op_protocol_data_4),
	.datab(avl_csr_address_2),
	.datac(\Selector27~4_combout ),
	.datad(csr_rd_inst_data_4),
	.cin(gnd),
	.combout(\Selector27~5_combout ),
	.cout());
defparam \Selector27~5 .lut_mask = 16'hF838;
defparam \Selector27~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector27~6 (
	.dataa(avl_csr_address_1),
	.datab(\Selector27~3_combout ),
	.datac(avl_csr_address_3),
	.datad(\Selector27~5_combout ),
	.cin(gnd),
	.combout(\Selector27~6_combout ),
	.cout());
defparam \Selector27~6 .lut_mask = 16'hE5E0;
defparam \Selector27~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector27~7 (
	.dataa(csr_flash_cmd_wr_data_1_data_4),
	.datab(csr_flash_cmd_wr_data_0_data_4),
	.datac(avl_csr_address_0),
	.datad(avl_csr_address_2),
	.cin(gnd),
	.combout(\Selector27~7_combout ),
	.cout());
defparam \Selector27~7 .lut_mask = 16'h00AC;
defparam \Selector27~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector27~8 (
	.dataa(\Selector27~1_combout ),
	.datab(avl_csr_address_1),
	.datac(\Selector27~6_combout ),
	.datad(\Selector27~7_combout ),
	.cin(gnd),
	.combout(\Selector27~8_combout ),
	.cout());
defparam \Selector27~8 .lut_mask = 16'hF838;
defparam \Selector27~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[4]~235 (
	.dataa(avl_csr_read),
	.datab(avl_csr_address_4),
	.datac(avl_csr_address_5),
	.datad(\Selector27~8_combout ),
	.cin(gnd),
	.combout(\rdata_comb[4]~235_combout ),
	.cout());
defparam \rdata_comb[4]~235 .lut_mask = 16'h0200;
defparam \rdata_comb[4]~235 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_csr_flash_cmd_addr~0 (
	.dataa(avl_csr_address_0),
	.datab(gnd),
	.datac(gnd),
	.datad(avl_csr_address_1),
	.cin(gnd),
	.combout(\wr_csr_flash_cmd_addr~0_combout ),
	.cout());
defparam \wr_csr_flash_cmd_addr~0 .lut_mask = 16'h00AA;
defparam \wr_csr_flash_cmd_addr~0 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[5] (
	.clk(clk),
	.d(out_rsp_data_5),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[5]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[5] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[5] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[5]~39 (
	.dataa(avl_csr_address_2),
	.datab(avl_csr_address_3),
	.datac(\wr_csr_flash_cmd_addr~0_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[5]~q ),
	.cin(gnd),
	.combout(\rdata_comb[5]~39_combout ),
	.cout());
defparam \rdata_comb[5]~39 .lut_mask = 16'h8000;
defparam \rdata_comb[5]~39 .sum_lutc_input = "datac";

cycloneive_lcell_comb \avl_rddata_local[7]~6 (
	.dataa(avl_csr_address_3),
	.datab(avl_csr_address_1),
	.datac(gnd),
	.datad(avl_csr_address_2),
	.cin(gnd),
	.combout(\avl_rddata_local[7]~6_combout ),
	.cout());
defparam \avl_rddata_local[7]~6 .lut_mask = 16'hAAEE;
defparam \avl_rddata_local[7]~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[5]~40 (
	.dataa(avl_csr_address_1),
	.datab(csr_rd_inst_data_5),
	.datac(avl_csr_address_0),
	.datad(csr_op_protocol_data_5),
	.cin(gnd),
	.combout(\rdata_comb[5]~40_combout ),
	.cout());
defparam \rdata_comb[5]~40 .lut_mask = 16'hE5E0;
defparam \rdata_comb[5]~40 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[5] (
	.clk(clk),
	.d(csr_wrdata[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[5]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[5] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[5] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[5]~41 (
	.dataa(csr_wr_inst_data_5),
	.datab(avl_csr_address_1),
	.datac(\rdata_comb[5]~40_combout ),
	.datad(\csr_flash_cmd_setting_data[5]~q ),
	.cin(gnd),
	.combout(\rdata_comb[5]~41_combout ),
	.cout());
defparam \rdata_comb[5]~41 .lut_mask = 16'hF838;
defparam \rdata_comb[5]~41 .sum_lutc_input = "datac";

cycloneive_lcell_comb \avl_rddata_local[7]~7 (
	.dataa(avl_csr_address_2),
	.datab(avl_csr_address_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\avl_rddata_local[7]~7_combout ),
	.cout());
defparam \avl_rddata_local[7]~7 .lut_mask = 16'hEEEE;
defparam \avl_rddata_local[7]~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[5]~42 (
	.dataa(\avl_rddata_local[7]~6_combout ),
	.datab(\rdata_comb[5]~41_combout ),
	.datac(\avl_rddata_local[7]~7_combout ),
	.datad(csr_control_data_5),
	.cin(gnd),
	.combout(\rdata_comb[5]~42_combout ),
	.cout());
defparam \rdata_comb[5]~42 .lut_mask = 16'hE5E0;
defparam \rdata_comb[5]~42 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_0_data[5] (
	.clk(clk),
	.d(out_rsp_data_5),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[5]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[5] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[5] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[5]~43 (
	.dataa(avl_csr_address_0),
	.datab(csr_flash_cmd_addr_data_5),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdata_comb[5]~43_combout ),
	.cout());
defparam \rdata_comb[5]~43 .lut_mask = 16'h8888;
defparam \rdata_comb[5]~43 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[5]~44 (
	.dataa(\csr_flash_cmd_rd_data_0_data[5]~q ),
	.datab(\rdata_comb[5]~43_combout ),
	.datac(avl_csr_address_1),
	.datad(\avl_rddata_local[3]~4_combout ),
	.cin(gnd),
	.combout(\rdata_comb[5]~44_combout ),
	.cout());
defparam \rdata_comb[5]~44 .lut_mask = 16'h0AFC;
defparam \rdata_comb[5]~44 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[5]~45 (
	.dataa(csr_flash_cmd_wr_data_1_data_5),
	.datab(csr_flash_cmd_wr_data_0_data_5),
	.datac(\avl_rddata_local[3]~3_combout ),
	.datad(\rdata_comb[5]~44_combout ),
	.cin(gnd),
	.combout(\rdata_comb[5]~45_combout ),
	.cout());
defparam \rdata_comb[5]~45 .lut_mask = 16'hCFA0;
defparam \rdata_comb[5]~45 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[5]~46 (
	.dataa(csr_delay_setting_data_5),
	.datab(\avl_rddata_local[7]~6_combout ),
	.datac(\rdata_comb[5]~42_combout ),
	.datad(\rdata_comb[5]~45_combout ),
	.cin(gnd),
	.combout(\rdata_comb[5]~46_combout ),
	.cout());
defparam \rdata_comb[5]~46 .lut_mask = 16'hF838;
defparam \rdata_comb[5]~46 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[5]~47 (
	.dataa(avl_csr_address_1),
	.datab(avl_csr_address_2),
	.datac(avl_csr_address_3),
	.datad(avl_csr_address_0),
	.cin(gnd),
	.combout(\rdata_comb[5]~47_combout ),
	.cout());
defparam \rdata_comb[5]~47 .lut_mask = 16'hBCFF;
defparam \rdata_comb[5]~47 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[5]~48 (
	.dataa(\rdata_comb[4]~10_combout ),
	.datab(\rdata_comb[5]~39_combout ),
	.datac(\rdata_comb[5]~46_combout ),
	.datad(\rdata_comb[5]~47_combout ),
	.cin(gnd),
	.combout(\rdata_comb[5]~48_combout ),
	.cout());
defparam \rdata_comb[5]~48 .lut_mask = 16'hA888;
defparam \rdata_comb[5]~48 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[6] (
	.clk(clk),
	.d(out_rsp_data_6),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[6]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[6] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[6] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[6]~49 (
	.dataa(avl_csr_address_2),
	.datab(avl_csr_address_3),
	.datac(\wr_csr_flash_cmd_addr~0_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[6]~q ),
	.cin(gnd),
	.combout(\rdata_comb[6]~49_combout ),
	.cout());
defparam \rdata_comb[6]~49 .lut_mask = 16'h8000;
defparam \rdata_comb[6]~49 .sum_lutc_input = "datac";

dffeas \csr_op_protocol_data[6] (
	.clk(clk),
	.d(csr_wrdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(\csr_op_protocol_data[6]~q ),
	.prn(vcc));
defparam \csr_op_protocol_data[6] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[6] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[6]~50 (
	.dataa(avl_csr_address_1),
	.datab(csr_rd_inst_data_6),
	.datac(avl_csr_address_0),
	.datad(\csr_op_protocol_data[6]~q ),
	.cin(gnd),
	.combout(\rdata_comb[6]~50_combout ),
	.cout());
defparam \rdata_comb[6]~50 .lut_mask = 16'hE5E0;
defparam \rdata_comb[6]~50 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[6] (
	.clk(clk),
	.d(csr_wrdata[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[6]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[6] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[6] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[6]~51 (
	.dataa(csr_wr_inst_data_6),
	.datab(avl_csr_address_1),
	.datac(\rdata_comb[6]~50_combout ),
	.datad(\csr_flash_cmd_setting_data[6]~q ),
	.cin(gnd),
	.combout(\rdata_comb[6]~51_combout ),
	.cout());
defparam \rdata_comb[6]~51 .lut_mask = 16'hF838;
defparam \rdata_comb[6]~51 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[6]~52 (
	.dataa(\avl_rddata_local[7]~7_combout ),
	.datab(csr_delay_setting_data_6),
	.datac(\avl_rddata_local[7]~6_combout ),
	.datad(csr_control_data_6),
	.cin(gnd),
	.combout(\rdata_comb[6]~52_combout ),
	.cout());
defparam \rdata_comb[6]~52 .lut_mask = 16'hE5E0;
defparam \rdata_comb[6]~52 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_0_data[6] (
	.clk(clk),
	.d(out_rsp_data_6),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[6]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[6] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[6] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[6]~53 (
	.dataa(avl_csr_address_0),
	.datab(csr_flash_cmd_addr_data_6),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdata_comb[6]~53_combout ),
	.cout());
defparam \rdata_comb[6]~53 .lut_mask = 16'h8888;
defparam \rdata_comb[6]~53 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[6]~54 (
	.dataa(\csr_flash_cmd_rd_data_0_data[6]~q ),
	.datab(\rdata_comb[6]~53_combout ),
	.datac(avl_csr_address_1),
	.datad(\avl_rddata_local[3]~4_combout ),
	.cin(gnd),
	.combout(\rdata_comb[6]~54_combout ),
	.cout());
defparam \rdata_comb[6]~54 .lut_mask = 16'h0AFC;
defparam \rdata_comb[6]~54 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[6]~55 (
	.dataa(csr_flash_cmd_wr_data_1_data_6),
	.datab(csr_flash_cmd_wr_data_0_data_6),
	.datac(\avl_rddata_local[3]~3_combout ),
	.datad(\rdata_comb[6]~54_combout ),
	.cin(gnd),
	.combout(\rdata_comb[6]~55_combout ),
	.cout());
defparam \rdata_comb[6]~55 .lut_mask = 16'hCFA0;
defparam \rdata_comb[6]~55 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[6]~56 (
	.dataa(\rdata_comb[6]~51_combout ),
	.datab(\avl_rddata_local[7]~7_combout ),
	.datac(\rdata_comb[6]~52_combout ),
	.datad(\rdata_comb[6]~55_combout ),
	.cin(gnd),
	.combout(\rdata_comb[6]~56_combout ),
	.cout());
defparam \rdata_comb[6]~56 .lut_mask = 16'hF838;
defparam \rdata_comb[6]~56 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[6]~57 (
	.dataa(\rdata_comb[4]~10_combout ),
	.datab(\rdata_comb[6]~49_combout ),
	.datac(\rdata_comb[5]~47_combout ),
	.datad(\rdata_comb[6]~56_combout ),
	.cin(gnd),
	.combout(\rdata_comb[6]~57_combout ),
	.cout());
defparam \rdata_comb[6]~57 .lut_mask = 16'hA888;
defparam \rdata_comb[6]~57 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[7] (
	.clk(clk),
	.d(out_rsp_data_7),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[7]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[7] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[7] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[7]~58 (
	.dataa(avl_csr_address_2),
	.datab(avl_csr_address_3),
	.datac(\wr_csr_flash_cmd_addr~0_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[7]~q ),
	.cin(gnd),
	.combout(\rdata_comb[7]~58_combout ),
	.cout());
defparam \rdata_comb[7]~58 .lut_mask = 16'h8000;
defparam \rdata_comb[7]~58 .sum_lutc_input = "datac";

dffeas \csr_op_protocol_data[7] (
	.clk(clk),
	.d(csr_wrdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(\csr_op_protocol_data[7]~q ),
	.prn(vcc));
defparam \csr_op_protocol_data[7] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[7] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[7]~59 (
	.dataa(avl_csr_address_1),
	.datab(csr_rd_inst_data_7),
	.datac(avl_csr_address_0),
	.datad(\csr_op_protocol_data[7]~q ),
	.cin(gnd),
	.combout(\rdata_comb[7]~59_combout ),
	.cout());
defparam \rdata_comb[7]~59 .lut_mask = 16'hE5E0;
defparam \rdata_comb[7]~59 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[7] (
	.clk(clk),
	.d(csr_wrdata[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[7]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[7] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[7] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[7]~60 (
	.dataa(csr_wr_inst_data_7),
	.datab(avl_csr_address_1),
	.datac(\rdata_comb[7]~59_combout ),
	.datad(\csr_flash_cmd_setting_data[7]~q ),
	.cin(gnd),
	.combout(\rdata_comb[7]~60_combout ),
	.cout());
defparam \rdata_comb[7]~60 .lut_mask = 16'hF838;
defparam \rdata_comb[7]~60 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[7]~61 (
	.dataa(\avl_rddata_local[7]~6_combout ),
	.datab(\rdata_comb[7]~60_combout ),
	.datac(\avl_rddata_local[7]~7_combout ),
	.datad(csr_control_data_7),
	.cin(gnd),
	.combout(\rdata_comb[7]~61_combout ),
	.cout());
defparam \rdata_comb[7]~61 .lut_mask = 16'hE5E0;
defparam \rdata_comb[7]~61 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_0_data[7] (
	.clk(clk),
	.d(out_rsp_data_7),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[7]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[7] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[7] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[7]~62 (
	.dataa(avl_csr_address_0),
	.datab(csr_flash_cmd_addr_data_7),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdata_comb[7]~62_combout ),
	.cout());
defparam \rdata_comb[7]~62 .lut_mask = 16'h8888;
defparam \rdata_comb[7]~62 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[7]~63 (
	.dataa(\csr_flash_cmd_rd_data_0_data[7]~q ),
	.datab(\rdata_comb[7]~62_combout ),
	.datac(avl_csr_address_1),
	.datad(\avl_rddata_local[3]~4_combout ),
	.cin(gnd),
	.combout(\rdata_comb[7]~63_combout ),
	.cout());
defparam \rdata_comb[7]~63 .lut_mask = 16'h0AFC;
defparam \rdata_comb[7]~63 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[7]~64 (
	.dataa(csr_flash_cmd_wr_data_1_data_7),
	.datab(csr_flash_cmd_wr_data_0_data_7),
	.datac(\avl_rddata_local[3]~3_combout ),
	.datad(\rdata_comb[7]~63_combout ),
	.cin(gnd),
	.combout(\rdata_comb[7]~64_combout ),
	.cout());
defparam \rdata_comb[7]~64 .lut_mask = 16'hCFA0;
defparam \rdata_comb[7]~64 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[7]~65 (
	.dataa(csr_delay_setting_data_7),
	.datab(\avl_rddata_local[7]~6_combout ),
	.datac(\rdata_comb[7]~61_combout ),
	.datad(\rdata_comb[7]~64_combout ),
	.cin(gnd),
	.combout(\rdata_comb[7]~65_combout ),
	.cout());
defparam \rdata_comb[7]~65 .lut_mask = 16'hF838;
defparam \rdata_comb[7]~65 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[7]~66 (
	.dataa(\rdata_comb[4]~10_combout ),
	.datab(\rdata_comb[7]~58_combout ),
	.datac(\rdata_comb[5]~47_combout ),
	.datad(\rdata_comb[7]~65_combout ),
	.cin(gnd),
	.combout(\rdata_comb[7]~66_combout ),
	.cout());
defparam \rdata_comb[7]~66 .lut_mask = 16'hA888;
defparam \rdata_comb[7]~66 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_0_data[8] (
	.clk(clk),
	.d(out_rsp_data_8),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[8]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[8] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[8] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[8]~67 (
	.dataa(avl_csr_address_3),
	.datab(csr_rd_inst_data_8),
	.datac(avl_csr_address_0),
	.datad(csr_op_protocol_data_8),
	.cin(gnd),
	.combout(\rdata_comb[8]~67_combout ),
	.cout());
defparam \rdata_comb[8]~67 .lut_mask = 16'hE5E0;
defparam \rdata_comb[8]~67 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[8] (
	.clk(clk),
	.d(out_rsp_data_8),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[8]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[8] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[8] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[8]~68 (
	.dataa(\csr_flash_cmd_rd_data_0_data[8]~q ),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[8]~67_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[8]~q ),
	.cin(gnd),
	.combout(\rdata_comb[8]~68_combout ),
	.cout());
defparam \rdata_comb[8]~68 .lut_mask = 16'hF838;
defparam \rdata_comb[8]~68 .sum_lutc_input = "datac";

cycloneive_lcell_comb \avl_rddata_local[13]~8 (
	.dataa(avl_csr_address_1),
	.datab(avl_csr_address_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\avl_rddata_local[13]~8_combout ),
	.cout());
defparam \avl_rddata_local[13]~8 .lut_mask = 16'hEEEE;
defparam \avl_rddata_local[13]~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \avl_rddata_local[13]~9 (
	.dataa(avl_csr_address_1),
	.datab(avl_csr_address_3),
	.datac(gnd),
	.datad(avl_csr_address_2),
	.cin(gnd),
	.combout(\avl_rddata_local[13]~9_combout ),
	.cout());
defparam \avl_rddata_local[13]~9 .lut_mask = 16'hAAEE;
defparam \avl_rddata_local[13]~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[8]~69 (
	.dataa(\avl_rddata_local[13]~8_combout ),
	.datab(csr_flash_cmd_addr_data_8),
	.datac(\avl_rddata_local[13]~9_combout ),
	.datad(csr_control_data_8),
	.cin(gnd),
	.combout(\rdata_comb[8]~69_combout ),
	.cout());
defparam \rdata_comb[8]~69 .lut_mask = 16'hE5E0;
defparam \rdata_comb[8]~69 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[8] (
	.clk(clk),
	.d(csr_wrdata[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[8]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[8] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[8] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[8]~70 (
	.dataa(avl_csr_address_3),
	.datab(\csr_flash_cmd_setting_data[8]~q ),
	.datac(avl_csr_address_0),
	.datad(csr_wr_inst_data_8),
	.cin(gnd),
	.combout(\rdata_comb[8]~70_combout ),
	.cout());
defparam \rdata_comb[8]~70 .lut_mask = 16'hE5E0;
defparam \rdata_comb[8]~70 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[8]~71 (
	.dataa(csr_flash_cmd_wr_data_0_data_8),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[8]~70_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_8),
	.cin(gnd),
	.combout(\rdata_comb[8]~71_combout ),
	.cout());
defparam \rdata_comb[8]~71 .lut_mask = 16'hF838;
defparam \rdata_comb[8]~71 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[8]~72 (
	.dataa(\rdata_comb[8]~68_combout ),
	.datab(\avl_rddata_local[13]~8_combout ),
	.datac(\rdata_comb[8]~69_combout ),
	.datad(\rdata_comb[8]~71_combout ),
	.cin(gnd),
	.combout(\rdata_comb[8]~72_combout ),
	.cout());
defparam \rdata_comb[8]~72 .lut_mask = 16'hF838;
defparam \rdata_comb[8]~72 .sum_lutc_input = "datac";

cycloneive_lcell_comb \avl_rddata_local[13]~11 (
	.dataa(avl_csr_address_1),
	.datab(avl_csr_address_3),
	.datac(avl_csr_address_2),
	.datad(avl_csr_address_0),
	.cin(gnd),
	.combout(\avl_rddata_local[13]~11_combout ),
	.cout());
defparam \avl_rddata_local[13]~11 .lut_mask = 16'hD9CC;
defparam \avl_rddata_local[13]~11 .sum_lutc_input = "datac";

cycloneive_lcell_comb \avl_rddata_local[13]~10 (
	.dataa(avl_csr_address_2),
	.datab(\rdata_comb[4]~10_combout ),
	.datac(avl_csr_address_1),
	.datad(\avl_rddata_local[13]~11_combout ),
	.cin(gnd),
	.combout(\avl_rddata_local[13]~10_combout ),
	.cout());
defparam \avl_rddata_local[13]~10 .lut_mask = 16'hB773;
defparam \avl_rddata_local[13]~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[8]~73 (
	.dataa(\rdata_comb[8]~72_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avl_rddata_local[13]~10_combout ),
	.cin(gnd),
	.combout(\rdata_comb[8]~73_combout ),
	.cout());
defparam \rdata_comb[8]~73 .lut_mask = 16'h00AA;
defparam \rdata_comb[8]~73 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_0_data[9] (
	.clk(clk),
	.d(out_rsp_data_9),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[9]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[9] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[9] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[9]~74 (
	.dataa(avl_csr_address_3),
	.datab(csr_rd_inst_data_9),
	.datac(avl_csr_address_0),
	.datad(csr_op_protocol_data_9),
	.cin(gnd),
	.combout(\rdata_comb[9]~74_combout ),
	.cout());
defparam \rdata_comb[9]~74 .lut_mask = 16'hE5E0;
defparam \rdata_comb[9]~74 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[9] (
	.clk(clk),
	.d(out_rsp_data_9),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[9]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[9] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[9] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[9]~75 (
	.dataa(\csr_flash_cmd_rd_data_0_data[9]~q ),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[9]~74_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[9]~q ),
	.cin(gnd),
	.combout(\rdata_comb[9]~75_combout ),
	.cout());
defparam \rdata_comb[9]~75 .lut_mask = 16'hF838;
defparam \rdata_comb[9]~75 .sum_lutc_input = "datac";

dffeas \csr_control_data[9] (
	.clk(clk),
	.d(csr_wrdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[9]~q ),
	.prn(vcc));
defparam \csr_control_data[9] .is_wysiwyg = "true";
defparam \csr_control_data[9] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[9]~76 (
	.dataa(\avl_rddata_local[13]~9_combout ),
	.datab(\rdata_comb[9]~75_combout ),
	.datac(\avl_rddata_local[13]~8_combout ),
	.datad(\csr_control_data[9]~q ),
	.cin(gnd),
	.combout(\rdata_comb[9]~76_combout ),
	.cout());
defparam \rdata_comb[9]~76 .lut_mask = 16'hE5E0;
defparam \rdata_comb[9]~76 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[9] (
	.clk(clk),
	.d(csr_wrdata[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[9]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[9] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[9] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[9]~77 (
	.dataa(avl_csr_address_3),
	.datab(\csr_flash_cmd_setting_data[9]~q ),
	.datac(avl_csr_address_0),
	.datad(csr_wr_inst_data_9),
	.cin(gnd),
	.combout(\rdata_comb[9]~77_combout ),
	.cout());
defparam \rdata_comb[9]~77 .lut_mask = 16'hE5E0;
defparam \rdata_comb[9]~77 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[9]~78 (
	.dataa(csr_flash_cmd_wr_data_0_data_9),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[9]~77_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_9),
	.cin(gnd),
	.combout(\rdata_comb[9]~78_combout ),
	.cout());
defparam \rdata_comb[9]~78 .lut_mask = 16'hF838;
defparam \rdata_comb[9]~78 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[9]~79 (
	.dataa(csr_flash_cmd_addr_data_9),
	.datab(\avl_rddata_local[13]~9_combout ),
	.datac(\rdata_comb[9]~76_combout ),
	.datad(\rdata_comb[9]~78_combout ),
	.cin(gnd),
	.combout(\rdata_comb[9]~79_combout ),
	.cout());
defparam \rdata_comb[9]~79 .lut_mask = 16'hF838;
defparam \rdata_comb[9]~79 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[9]~80 (
	.dataa(\rdata_comb[9]~79_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avl_rddata_local[13]~10_combout ),
	.cin(gnd),
	.combout(\rdata_comb[9]~80_combout ),
	.cout());
defparam \rdata_comb[9]~80 .lut_mask = 16'h00AA;
defparam \rdata_comb[9]~80 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_0_data[10] (
	.clk(clk),
	.d(out_rsp_data_10),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[10]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[10] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[10] .power_up = "low";

dffeas \csr_op_protocol_data[10] (
	.clk(clk),
	.d(csr_wrdata[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(\csr_op_protocol_data[10]~q ),
	.prn(vcc));
defparam \csr_op_protocol_data[10] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[10] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[10]~81 (
	.dataa(avl_csr_address_3),
	.datab(csr_rd_inst_data_10),
	.datac(avl_csr_address_0),
	.datad(\csr_op_protocol_data[10]~q ),
	.cin(gnd),
	.combout(\rdata_comb[10]~81_combout ),
	.cout());
defparam \rdata_comb[10]~81 .lut_mask = 16'hE5E0;
defparam \rdata_comb[10]~81 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[10] (
	.clk(clk),
	.d(out_rsp_data_10),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[10]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[10] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[10] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[10]~82 (
	.dataa(\csr_flash_cmd_rd_data_0_data[10]~q ),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[10]~81_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[10]~q ),
	.cin(gnd),
	.combout(\rdata_comb[10]~82_combout ),
	.cout());
defparam \rdata_comb[10]~82 .lut_mask = 16'hF838;
defparam \rdata_comb[10]~82 .sum_lutc_input = "datac";

dffeas \csr_control_data[10] (
	.clk(clk),
	.d(csr_wrdata[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[10]~q ),
	.prn(vcc));
defparam \csr_control_data[10] .is_wysiwyg = "true";
defparam \csr_control_data[10] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[10]~83 (
	.dataa(\avl_rddata_local[13]~8_combout ),
	.datab(csr_flash_cmd_addr_data_10),
	.datac(\avl_rddata_local[13]~9_combout ),
	.datad(\csr_control_data[10]~q ),
	.cin(gnd),
	.combout(\rdata_comb[10]~83_combout ),
	.cout());
defparam \rdata_comb[10]~83 .lut_mask = 16'hE5E0;
defparam \rdata_comb[10]~83 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[10] (
	.clk(clk),
	.d(csr_wrdata[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[10]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[10] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[10] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[10]~84 (
	.dataa(avl_csr_address_3),
	.datab(\csr_flash_cmd_setting_data[10]~q ),
	.datac(avl_csr_address_0),
	.datad(csr_wr_inst_data_10),
	.cin(gnd),
	.combout(\rdata_comb[10]~84_combout ),
	.cout());
defparam \rdata_comb[10]~84 .lut_mask = 16'hE5E0;
defparam \rdata_comb[10]~84 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[10]~85 (
	.dataa(csr_flash_cmd_wr_data_0_data_10),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[10]~84_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_10),
	.cin(gnd),
	.combout(\rdata_comb[10]~85_combout ),
	.cout());
defparam \rdata_comb[10]~85 .lut_mask = 16'hF838;
defparam \rdata_comb[10]~85 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[10]~86 (
	.dataa(\rdata_comb[10]~82_combout ),
	.datab(\avl_rddata_local[13]~8_combout ),
	.datac(\rdata_comb[10]~83_combout ),
	.datad(\rdata_comb[10]~85_combout ),
	.cin(gnd),
	.combout(\rdata_comb[10]~86_combout ),
	.cout());
defparam \rdata_comb[10]~86 .lut_mask = 16'hF838;
defparam \rdata_comb[10]~86 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[10]~87 (
	.dataa(\rdata_comb[10]~86_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avl_rddata_local[13]~10_combout ),
	.cin(gnd),
	.combout(\rdata_comb[10]~87_combout ),
	.cout());
defparam \rdata_comb[10]~87 .lut_mask = 16'h00AA;
defparam \rdata_comb[10]~87 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_0_data[11] (
	.clk(clk),
	.d(out_rsp_data_11),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[11]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[11] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[11] .power_up = "low";

dffeas \csr_op_protocol_data[11] (
	.clk(clk),
	.d(csr_wrdata[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(\csr_op_protocol_data[11]~q ),
	.prn(vcc));
defparam \csr_op_protocol_data[11] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[11] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[11]~88 (
	.dataa(avl_csr_address_3),
	.datab(csr_rd_inst_data_11),
	.datac(avl_csr_address_0),
	.datad(\csr_op_protocol_data[11]~q ),
	.cin(gnd),
	.combout(\rdata_comb[11]~88_combout ),
	.cout());
defparam \rdata_comb[11]~88 .lut_mask = 16'hE5E0;
defparam \rdata_comb[11]~88 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[11] (
	.clk(clk),
	.d(out_rsp_data_11),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[11]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[11] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[11] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[11]~89 (
	.dataa(\csr_flash_cmd_rd_data_0_data[11]~q ),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[11]~88_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[11]~q ),
	.cin(gnd),
	.combout(\rdata_comb[11]~89_combout ),
	.cout());
defparam \rdata_comb[11]~89 .lut_mask = 16'hF838;
defparam \rdata_comb[11]~89 .sum_lutc_input = "datac";

dffeas \csr_control_data[11] (
	.clk(clk),
	.d(csr_wrdata[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[11]~q ),
	.prn(vcc));
defparam \csr_control_data[11] .is_wysiwyg = "true";
defparam \csr_control_data[11] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[11]~90 (
	.dataa(\avl_rddata_local[13]~9_combout ),
	.datab(\rdata_comb[11]~89_combout ),
	.datac(\avl_rddata_local[13]~8_combout ),
	.datad(\csr_control_data[11]~q ),
	.cin(gnd),
	.combout(\rdata_comb[11]~90_combout ),
	.cout());
defparam \rdata_comb[11]~90 .lut_mask = 16'hE5E0;
defparam \rdata_comb[11]~90 .sum_lutc_input = "datac";

cycloneive_lcell_comb \csr_flash_cmd_setting_data[11]~2 (
	.dataa(csr_wrdata[11]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\csr_flash_cmd_setting_data[11]~2_combout ),
	.cout());
defparam \csr_flash_cmd_setting_data[11]~2 .lut_mask = 16'h5555;
defparam \csr_flash_cmd_setting_data[11]~2 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[11] (
	.clk(clk),
	.d(\csr_flash_cmd_setting_data[11]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[11]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[11] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[11] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[11]~91 (
	.dataa(avl_csr_address_3),
	.datab(\csr_flash_cmd_setting_data[11]~q ),
	.datac(avl_csr_address_0),
	.datad(csr_wr_inst_data_11),
	.cin(gnd),
	.combout(\rdata_comb[11]~91_combout ),
	.cout());
defparam \rdata_comb[11]~91 .lut_mask = 16'hB5B0;
defparam \rdata_comb[11]~91 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[11]~92 (
	.dataa(csr_flash_cmd_wr_data_0_data_11),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[11]~91_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_11),
	.cin(gnd),
	.combout(\rdata_comb[11]~92_combout ),
	.cout());
defparam \rdata_comb[11]~92 .lut_mask = 16'hF838;
defparam \rdata_comb[11]~92 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[11]~93 (
	.dataa(csr_flash_cmd_addr_data_11),
	.datab(\avl_rddata_local[13]~9_combout ),
	.datac(\rdata_comb[11]~90_combout ),
	.datad(\rdata_comb[11]~92_combout ),
	.cin(gnd),
	.combout(\rdata_comb[11]~93_combout ),
	.cout());
defparam \rdata_comb[11]~93 .lut_mask = 16'hF838;
defparam \rdata_comb[11]~93 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[11]~94 (
	.dataa(\rdata_comb[11]~93_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avl_rddata_local[13]~10_combout ),
	.cin(gnd),
	.combout(\rdata_comb[11]~94_combout ),
	.cout());
defparam \rdata_comb[11]~94 .lut_mask = 16'h00AA;
defparam \rdata_comb[11]~94 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_0_data[12] (
	.clk(clk),
	.d(out_rsp_data_12),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[12]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[12] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[12] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[12]~95 (
	.dataa(avl_csr_address_3),
	.datab(csr_rd_inst_data_12),
	.datac(avl_csr_address_0),
	.datad(csr_op_protocol_data_12),
	.cin(gnd),
	.combout(\rdata_comb[12]~95_combout ),
	.cout());
defparam \rdata_comb[12]~95 .lut_mask = 16'hE5E0;
defparam \rdata_comb[12]~95 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[12] (
	.clk(clk),
	.d(out_rsp_data_12),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[12]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[12] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[12] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[12]~96 (
	.dataa(\csr_flash_cmd_rd_data_0_data[12]~q ),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[12]~95_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[12]~q ),
	.cin(gnd),
	.combout(\rdata_comb[12]~96_combout ),
	.cout());
defparam \rdata_comb[12]~96 .lut_mask = 16'hF838;
defparam \rdata_comb[12]~96 .sum_lutc_input = "datac";

dffeas \csr_control_data[12] (
	.clk(clk),
	.d(csr_wrdata[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[12]~q ),
	.prn(vcc));
defparam \csr_control_data[12] .is_wysiwyg = "true";
defparam \csr_control_data[12] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[12]~97 (
	.dataa(\avl_rddata_local[13]~8_combout ),
	.datab(csr_flash_cmd_addr_data_12),
	.datac(\avl_rddata_local[13]~9_combout ),
	.datad(\csr_control_data[12]~q ),
	.cin(gnd),
	.combout(\rdata_comb[12]~97_combout ),
	.cout());
defparam \rdata_comb[12]~97 .lut_mask = 16'hE5E0;
defparam \rdata_comb[12]~97 .sum_lutc_input = "datac";

cycloneive_lcell_comb \csr_flash_cmd_setting_data[12]~3 (
	.dataa(csr_wrdata[12]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\csr_flash_cmd_setting_data[12]~3_combout ),
	.cout());
defparam \csr_flash_cmd_setting_data[12]~3 .lut_mask = 16'h5555;
defparam \csr_flash_cmd_setting_data[12]~3 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[12] (
	.clk(clk),
	.d(\csr_flash_cmd_setting_data[12]~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[12]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[12] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[12] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[12]~98 (
	.dataa(avl_csr_address_3),
	.datab(\csr_flash_cmd_setting_data[12]~q ),
	.datac(avl_csr_address_0),
	.datad(csr_wr_inst_data_12),
	.cin(gnd),
	.combout(\rdata_comb[12]~98_combout ),
	.cout());
defparam \rdata_comb[12]~98 .lut_mask = 16'hB0B5;
defparam \rdata_comb[12]~98 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[12]~99 (
	.dataa(csr_flash_cmd_wr_data_0_data_12),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[12]~98_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_12),
	.cin(gnd),
	.combout(\rdata_comb[12]~99_combout ),
	.cout());
defparam \rdata_comb[12]~99 .lut_mask = 16'hF838;
defparam \rdata_comb[12]~99 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[12]~100 (
	.dataa(\rdata_comb[12]~96_combout ),
	.datab(\avl_rddata_local[13]~8_combout ),
	.datac(\rdata_comb[12]~97_combout ),
	.datad(\rdata_comb[12]~99_combout ),
	.cin(gnd),
	.combout(\rdata_comb[12]~100_combout ),
	.cout());
defparam \rdata_comb[12]~100 .lut_mask = 16'hF838;
defparam \rdata_comb[12]~100 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[12]~101 (
	.dataa(\rdata_comb[12]~100_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avl_rddata_local[13]~10_combout ),
	.cin(gnd),
	.combout(\rdata_comb[12]~101_combout ),
	.cout());
defparam \rdata_comb[12]~101 .lut_mask = 16'h00AA;
defparam \rdata_comb[12]~101 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_0_data[13] (
	.clk(clk),
	.d(out_rsp_data_13),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[13]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[13] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[13] .power_up = "low";

cycloneive_lcell_comb wr_csr_rd_inst(
	.dataa(avl_csr_address_2),
	.datab(\wr_csr_flash_cmd_addr~0_combout ),
	.datac(\wr_csr_control~0_combout ),
	.datad(avl_csr_address_3),
	.cin(gnd),
	.combout(\wr_csr_rd_inst~combout ),
	.cout());
defparam wr_csr_rd_inst.lut_mask = 16'h0080;
defparam wr_csr_rd_inst.sum_lutc_input = "datac";

dffeas \csr_rd_inst_data[13] (
	.clk(clk),
	.d(csr_wrdata[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(\csr_rd_inst_data[13]~q ),
	.prn(vcc));
defparam \csr_rd_inst_data[13] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[13] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[13]~102 (
	.dataa(avl_csr_address_3),
	.datab(\csr_rd_inst_data[13]~q ),
	.datac(avl_csr_address_0),
	.datad(csr_op_protocol_data_13),
	.cin(gnd),
	.combout(\rdata_comb[13]~102_combout ),
	.cout());
defparam \rdata_comb[13]~102 .lut_mask = 16'hE5E0;
defparam \rdata_comb[13]~102 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[13] (
	.clk(clk),
	.d(out_rsp_data_13),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[13]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[13] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[13] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[13]~103 (
	.dataa(\csr_flash_cmd_rd_data_0_data[13]~q ),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[13]~102_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[13]~q ),
	.cin(gnd),
	.combout(\rdata_comb[13]~103_combout ),
	.cout());
defparam \rdata_comb[13]~103 .lut_mask = 16'hF838;
defparam \rdata_comb[13]~103 .sum_lutc_input = "datac";

dffeas \csr_control_data[13] (
	.clk(clk),
	.d(csr_wrdata[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[13]~q ),
	.prn(vcc));
defparam \csr_control_data[13] .is_wysiwyg = "true";
defparam \csr_control_data[13] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[13]~104 (
	.dataa(\avl_rddata_local[13]~9_combout ),
	.datab(\rdata_comb[13]~103_combout ),
	.datac(\avl_rddata_local[13]~8_combout ),
	.datad(\csr_control_data[13]~q ),
	.cin(gnd),
	.combout(\rdata_comb[13]~104_combout ),
	.cout());
defparam \rdata_comb[13]~104 .lut_mask = 16'hE5E0;
defparam \rdata_comb[13]~104 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[13] (
	.clk(clk),
	.d(csr_wrdata[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[13]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[13] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[13] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[13]~105 (
	.dataa(avl_csr_address_3),
	.datab(\csr_flash_cmd_setting_data[13]~q ),
	.datac(avl_csr_address_0),
	.datad(csr_wr_inst_data_13),
	.cin(gnd),
	.combout(\rdata_comb[13]~105_combout ),
	.cout());
defparam \rdata_comb[13]~105 .lut_mask = 16'hE0E5;
defparam \rdata_comb[13]~105 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[13]~106 (
	.dataa(csr_flash_cmd_wr_data_0_data_13),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[13]~105_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_13),
	.cin(gnd),
	.combout(\rdata_comb[13]~106_combout ),
	.cout());
defparam \rdata_comb[13]~106 .lut_mask = 16'hF838;
defparam \rdata_comb[13]~106 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[13]~107 (
	.dataa(csr_flash_cmd_addr_data_13),
	.datab(\avl_rddata_local[13]~9_combout ),
	.datac(\rdata_comb[13]~104_combout ),
	.datad(\rdata_comb[13]~106_combout ),
	.cin(gnd),
	.combout(\rdata_comb[13]~107_combout ),
	.cout());
defparam \rdata_comb[13]~107 .lut_mask = 16'hF838;
defparam \rdata_comb[13]~107 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[13]~108 (
	.dataa(\rdata_comb[13]~107_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avl_rddata_local[13]~10_combout ),
	.cin(gnd),
	.combout(\rdata_comb[13]~108_combout ),
	.cout());
defparam \rdata_comb[13]~108 .lut_mask = 16'h00AA;
defparam \rdata_comb[13]~108 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_0_data[14] (
	.clk(clk),
	.d(out_rsp_data_14),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[14]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[14] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[14] .power_up = "low";

dffeas \csr_rd_inst_data[14] (
	.clk(clk),
	.d(csr_wrdata[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(\csr_rd_inst_data[14]~q ),
	.prn(vcc));
defparam \csr_rd_inst_data[14] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[14] .power_up = "low";

dffeas \csr_op_protocol_data[14] (
	.clk(clk),
	.d(csr_wrdata[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(\csr_op_protocol_data[14]~q ),
	.prn(vcc));
defparam \csr_op_protocol_data[14] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[14] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[14]~109 (
	.dataa(avl_csr_address_3),
	.datab(\csr_rd_inst_data[14]~q ),
	.datac(avl_csr_address_0),
	.datad(\csr_op_protocol_data[14]~q ),
	.cin(gnd),
	.combout(\rdata_comb[14]~109_combout ),
	.cout());
defparam \rdata_comb[14]~109 .lut_mask = 16'hE5E0;
defparam \rdata_comb[14]~109 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[14] (
	.clk(clk),
	.d(out_rsp_data_14),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[14]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[14] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[14] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[14]~110 (
	.dataa(\csr_flash_cmd_rd_data_0_data[14]~q ),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[14]~109_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[14]~q ),
	.cin(gnd),
	.combout(\rdata_comb[14]~110_combout ),
	.cout());
defparam \rdata_comb[14]~110 .lut_mask = 16'hF838;
defparam \rdata_comb[14]~110 .sum_lutc_input = "datac";

dffeas \csr_control_data[14] (
	.clk(clk),
	.d(csr_wrdata[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[14]~q ),
	.prn(vcc));
defparam \csr_control_data[14] .is_wysiwyg = "true";
defparam \csr_control_data[14] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[14]~111 (
	.dataa(\avl_rddata_local[13]~8_combout ),
	.datab(csr_flash_cmd_addr_data_14),
	.datac(\avl_rddata_local[13]~9_combout ),
	.datad(\csr_control_data[14]~q ),
	.cin(gnd),
	.combout(\rdata_comb[14]~111_combout ),
	.cout());
defparam \rdata_comb[14]~111 .lut_mask = 16'hE5E0;
defparam \rdata_comb[14]~111 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[14] (
	.clk(clk),
	.d(csr_wrdata[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[14]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[14] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[14] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[14]~112 (
	.dataa(avl_csr_address_3),
	.datab(\csr_flash_cmd_setting_data[14]~q ),
	.datac(avl_csr_address_0),
	.datad(csr_wr_inst_data_14),
	.cin(gnd),
	.combout(\rdata_comb[14]~112_combout ),
	.cout());
defparam \rdata_comb[14]~112 .lut_mask = 16'hE0E5;
defparam \rdata_comb[14]~112 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[14]~113 (
	.dataa(csr_flash_cmd_wr_data_0_data_14),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[14]~112_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_14),
	.cin(gnd),
	.combout(\rdata_comb[14]~113_combout ),
	.cout());
defparam \rdata_comb[14]~113 .lut_mask = 16'hF838;
defparam \rdata_comb[14]~113 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[14]~114 (
	.dataa(\rdata_comb[14]~110_combout ),
	.datab(\avl_rddata_local[13]~8_combout ),
	.datac(\rdata_comb[14]~111_combout ),
	.datad(\rdata_comb[14]~113_combout ),
	.cin(gnd),
	.combout(\rdata_comb[14]~114_combout ),
	.cout());
defparam \rdata_comb[14]~114 .lut_mask = 16'hF838;
defparam \rdata_comb[14]~114 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[14]~115 (
	.dataa(\rdata_comb[14]~114_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avl_rddata_local[13]~10_combout ),
	.cin(gnd),
	.combout(\rdata_comb[14]~115_combout ),
	.cout());
defparam \rdata_comb[14]~115 .lut_mask = 16'h00AA;
defparam \rdata_comb[14]~115 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_0_data[15] (
	.clk(clk),
	.d(out_rsp_data_15),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[15]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[15] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[15] .power_up = "low";

dffeas \csr_rd_inst_data[15] (
	.clk(clk),
	.d(csr_wrdata[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(\csr_rd_inst_data[15]~q ),
	.prn(vcc));
defparam \csr_rd_inst_data[15] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[15] .power_up = "low";

dffeas \csr_op_protocol_data[15] (
	.clk(clk),
	.d(csr_wrdata[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(\csr_op_protocol_data[15]~q ),
	.prn(vcc));
defparam \csr_op_protocol_data[15] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[15] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[15]~116 (
	.dataa(avl_csr_address_3),
	.datab(\csr_rd_inst_data[15]~q ),
	.datac(avl_csr_address_0),
	.datad(\csr_op_protocol_data[15]~q ),
	.cin(gnd),
	.combout(\rdata_comb[15]~116_combout ),
	.cout());
defparam \rdata_comb[15]~116 .lut_mask = 16'hE5E0;
defparam \rdata_comb[15]~116 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[15] (
	.clk(clk),
	.d(out_rsp_data_15),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[15]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[15] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[15] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[15]~117 (
	.dataa(\csr_flash_cmd_rd_data_0_data[15]~q ),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[15]~116_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[15]~q ),
	.cin(gnd),
	.combout(\rdata_comb[15]~117_combout ),
	.cout());
defparam \rdata_comb[15]~117 .lut_mask = 16'hF838;
defparam \rdata_comb[15]~117 .sum_lutc_input = "datac";

dffeas \csr_control_data[15] (
	.clk(clk),
	.d(csr_wrdata[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[15]~q ),
	.prn(vcc));
defparam \csr_control_data[15] .is_wysiwyg = "true";
defparam \csr_control_data[15] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[15]~118 (
	.dataa(\avl_rddata_local[13]~9_combout ),
	.datab(\rdata_comb[15]~117_combout ),
	.datac(\avl_rddata_local[13]~8_combout ),
	.datad(\csr_control_data[15]~q ),
	.cin(gnd),
	.combout(\rdata_comb[15]~118_combout ),
	.cout());
defparam \rdata_comb[15]~118 .lut_mask = 16'hE5E0;
defparam \rdata_comb[15]~118 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[15] (
	.clk(clk),
	.d(csr_wrdata[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[15]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[15] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[15] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[15]~119 (
	.dataa(avl_csr_address_3),
	.datab(\csr_flash_cmd_setting_data[15]~q ),
	.datac(avl_csr_address_0),
	.datad(csr_wr_inst_data_15),
	.cin(gnd),
	.combout(\rdata_comb[15]~119_combout ),
	.cout());
defparam \rdata_comb[15]~119 .lut_mask = 16'hE5E0;
defparam \rdata_comb[15]~119 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[15]~120 (
	.dataa(csr_flash_cmd_wr_data_0_data_15),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[15]~119_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_15),
	.cin(gnd),
	.combout(\rdata_comb[15]~120_combout ),
	.cout());
defparam \rdata_comb[15]~120 .lut_mask = 16'hF838;
defparam \rdata_comb[15]~120 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[15]~121 (
	.dataa(csr_flash_cmd_addr_data_15),
	.datab(\avl_rddata_local[13]~9_combout ),
	.datac(\rdata_comb[15]~118_combout ),
	.datad(\rdata_comb[15]~120_combout ),
	.cin(gnd),
	.combout(\rdata_comb[15]~121_combout ),
	.cout());
defparam \rdata_comb[15]~121 .lut_mask = 16'hF838;
defparam \rdata_comb[15]~121 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[15]~122 (
	.dataa(\rdata_comb[15]~121_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avl_rddata_local[13]~10_combout ),
	.cin(gnd),
	.combout(\rdata_comb[15]~122_combout ),
	.cout());
defparam \rdata_comb[15]~122 .lut_mask = 16'h00AA;
defparam \rdata_comb[15]~122 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_0_data[16] (
	.clk(clk),
	.d(out_rsp_data_16),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[16]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[16] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[16] .power_up = "low";

dffeas \csr_rd_inst_data[16] (
	.clk(clk),
	.d(csr_wrdata[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(\csr_rd_inst_data[16]~q ),
	.prn(vcc));
defparam \csr_rd_inst_data[16] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[16] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[16]~123 (
	.dataa(avl_csr_address_3),
	.datab(\csr_rd_inst_data[16]~q ),
	.datac(avl_csr_address_0),
	.datad(csr_op_protocol_data_16),
	.cin(gnd),
	.combout(\rdata_comb[16]~123_combout ),
	.cout());
defparam \rdata_comb[16]~123 .lut_mask = 16'hE5E0;
defparam \rdata_comb[16]~123 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[16] (
	.clk(clk),
	.d(out_rsp_data_16),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[16]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[16] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[16] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[16]~124 (
	.dataa(\csr_flash_cmd_rd_data_0_data[16]~q ),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[16]~123_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[16]~q ),
	.cin(gnd),
	.combout(\rdata_comb[16]~124_combout ),
	.cout());
defparam \rdata_comb[16]~124 .lut_mask = 16'hF838;
defparam \rdata_comb[16]~124 .sum_lutc_input = "datac";

dffeas \csr_control_data[16] (
	.clk(clk),
	.d(csr_wrdata[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[16]~q ),
	.prn(vcc));
defparam \csr_control_data[16] .is_wysiwyg = "true";
defparam \csr_control_data[16] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[16]~125 (
	.dataa(\avl_rddata_local[13]~8_combout ),
	.datab(csr_flash_cmd_addr_data_16),
	.datac(\avl_rddata_local[13]~9_combout ),
	.datad(\csr_control_data[16]~q ),
	.cin(gnd),
	.combout(\rdata_comb[16]~125_combout ),
	.cout());
defparam \rdata_comb[16]~125 .lut_mask = 16'hE5E0;
defparam \rdata_comb[16]~125 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[16] (
	.clk(clk),
	.d(csr_wrdata[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[16]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[16] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[16] .power_up = "low";

cycloneive_lcell_comb wr_csr_wr_inst(
	.dataa(avl_csr_address_1),
	.datab(\wr_csr_op_protocol~0_combout ),
	.datac(gnd),
	.datad(avl_csr_address_0),
	.cin(gnd),
	.combout(\wr_csr_wr_inst~combout ),
	.cout());
defparam wr_csr_wr_inst.lut_mask = 16'h0088;
defparam wr_csr_wr_inst.sum_lutc_input = "datac";

dffeas \csr_wr_inst_data[16] (
	.clk(clk),
	.d(csr_wrdata[16]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(\csr_wr_inst_data[16]~q ),
	.prn(vcc));
defparam \csr_wr_inst_data[16] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[16] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[16]~126 (
	.dataa(avl_csr_address_3),
	.datab(\csr_flash_cmd_setting_data[16]~q ),
	.datac(avl_csr_address_0),
	.datad(\csr_wr_inst_data[16]~q ),
	.cin(gnd),
	.combout(\rdata_comb[16]~126_combout ),
	.cout());
defparam \rdata_comb[16]~126 .lut_mask = 16'hE5E0;
defparam \rdata_comb[16]~126 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[16]~127 (
	.dataa(csr_flash_cmd_wr_data_0_data_16),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[16]~126_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_16),
	.cin(gnd),
	.combout(\rdata_comb[16]~127_combout ),
	.cout());
defparam \rdata_comb[16]~127 .lut_mask = 16'hF838;
defparam \rdata_comb[16]~127 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[16]~128 (
	.dataa(\rdata_comb[16]~124_combout ),
	.datab(\avl_rddata_local[13]~8_combout ),
	.datac(\rdata_comb[16]~125_combout ),
	.datad(\rdata_comb[16]~127_combout ),
	.cin(gnd),
	.combout(\rdata_comb[16]~128_combout ),
	.cout());
defparam \rdata_comb[16]~128 .lut_mask = 16'hF838;
defparam \rdata_comb[16]~128 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[16]~129 (
	.dataa(\rdata_comb[16]~128_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avl_rddata_local[13]~10_combout ),
	.cin(gnd),
	.combout(\rdata_comb[16]~129_combout ),
	.cout());
defparam \rdata_comb[16]~129 .lut_mask = 16'h00AA;
defparam \rdata_comb[16]~129 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_0_data[17] (
	.clk(clk),
	.d(out_rsp_data_17),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[17]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[17] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[17] .power_up = "low";

dffeas \csr_rd_inst_data[17] (
	.clk(clk),
	.d(csr_wrdata[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(\csr_rd_inst_data[17]~q ),
	.prn(vcc));
defparam \csr_rd_inst_data[17] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[17] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[17]~130 (
	.dataa(avl_csr_address_3),
	.datab(\csr_rd_inst_data[17]~q ),
	.datac(avl_csr_address_0),
	.datad(csr_op_protocol_data_17),
	.cin(gnd),
	.combout(\rdata_comb[17]~130_combout ),
	.cout());
defparam \rdata_comb[17]~130 .lut_mask = 16'hE5E0;
defparam \rdata_comb[17]~130 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[17] (
	.clk(clk),
	.d(out_rsp_data_17),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[17]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[17] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[17] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[17]~131 (
	.dataa(\csr_flash_cmd_rd_data_0_data[17]~q ),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[17]~130_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[17]~q ),
	.cin(gnd),
	.combout(\rdata_comb[17]~131_combout ),
	.cout());
defparam \rdata_comb[17]~131 .lut_mask = 16'hF838;
defparam \rdata_comb[17]~131 .sum_lutc_input = "datac";

dffeas \csr_control_data[17] (
	.clk(clk),
	.d(csr_wrdata[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[17]~q ),
	.prn(vcc));
defparam \csr_control_data[17] .is_wysiwyg = "true";
defparam \csr_control_data[17] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[17]~132 (
	.dataa(\avl_rddata_local[13]~9_combout ),
	.datab(\rdata_comb[17]~131_combout ),
	.datac(\avl_rddata_local[13]~8_combout ),
	.datad(\csr_control_data[17]~q ),
	.cin(gnd),
	.combout(\rdata_comb[17]~132_combout ),
	.cout());
defparam \rdata_comb[17]~132 .lut_mask = 16'hE5E0;
defparam \rdata_comb[17]~132 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[17] (
	.clk(clk),
	.d(csr_wrdata[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[17]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[17] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[17] .power_up = "low";

dffeas \csr_wr_inst_data[17] (
	.clk(clk),
	.d(csr_wrdata[17]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(\csr_wr_inst_data[17]~q ),
	.prn(vcc));
defparam \csr_wr_inst_data[17] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[17] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[17]~133 (
	.dataa(avl_csr_address_3),
	.datab(\csr_flash_cmd_setting_data[17]~q ),
	.datac(avl_csr_address_0),
	.datad(\csr_wr_inst_data[17]~q ),
	.cin(gnd),
	.combout(\rdata_comb[17]~133_combout ),
	.cout());
defparam \rdata_comb[17]~133 .lut_mask = 16'hE5E0;
defparam \rdata_comb[17]~133 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[17]~134 (
	.dataa(csr_flash_cmd_wr_data_0_data_17),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[17]~133_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_17),
	.cin(gnd),
	.combout(\rdata_comb[17]~134_combout ),
	.cout());
defparam \rdata_comb[17]~134 .lut_mask = 16'hF838;
defparam \rdata_comb[17]~134 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[17]~135 (
	.dataa(csr_flash_cmd_addr_data_17),
	.datab(\avl_rddata_local[13]~9_combout ),
	.datac(\rdata_comb[17]~132_combout ),
	.datad(\rdata_comb[17]~134_combout ),
	.cin(gnd),
	.combout(\rdata_comb[17]~135_combout ),
	.cout());
defparam \rdata_comb[17]~135 .lut_mask = 16'hF838;
defparam \rdata_comb[17]~135 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[17]~136 (
	.dataa(\rdata_comb[17]~135_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avl_rddata_local[13]~10_combout ),
	.cin(gnd),
	.combout(\rdata_comb[17]~136_combout ),
	.cout());
defparam \rdata_comb[17]~136 .lut_mask = 16'h00AA;
defparam \rdata_comb[17]~136 .sum_lutc_input = "datac";

dffeas \csr_rd_inst_data[18] (
	.clk(clk),
	.d(csr_wrdata[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(\csr_rd_inst_data[18]~q ),
	.prn(vcc));
defparam \csr_rd_inst_data[18] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[18] .power_up = "low";

dffeas \csr_flash_cmd_rd_data_0_data[18] (
	.clk(clk),
	.d(out_rsp_data_18),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[18]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[18] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[18] .power_up = "low";

dffeas \csr_op_protocol_data[18] (
	.clk(clk),
	.d(csr_wrdata[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(\csr_op_protocol_data[18]~q ),
	.prn(vcc));
defparam \csr_op_protocol_data[18] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[18] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[18]~137 (
	.dataa(avl_csr_address_0),
	.datab(\csr_flash_cmd_rd_data_0_data[18]~q ),
	.datac(avl_csr_address_3),
	.datad(\csr_op_protocol_data[18]~q ),
	.cin(gnd),
	.combout(\rdata_comb[18]~137_combout ),
	.cout());
defparam \rdata_comb[18]~137 .lut_mask = 16'hE5E0;
defparam \rdata_comb[18]~137 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[18] (
	.clk(clk),
	.d(out_rsp_data_18),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[18]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[18] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[18] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[18]~138 (
	.dataa(\csr_rd_inst_data[18]~q ),
	.datab(avl_csr_address_0),
	.datac(\rdata_comb[18]~137_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[18]~q ),
	.cin(gnd),
	.combout(\rdata_comb[18]~138_combout ),
	.cout());
defparam \rdata_comb[18]~138 .lut_mask = 16'hF838;
defparam \rdata_comb[18]~138 .sum_lutc_input = "datac";

dffeas \csr_control_data[18] (
	.clk(clk),
	.d(csr_wrdata[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[18]~q ),
	.prn(vcc));
defparam \csr_control_data[18] .is_wysiwyg = "true";
defparam \csr_control_data[18] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[18]~139 (
	.dataa(\avl_rddata_local[13]~8_combout ),
	.datab(csr_flash_cmd_addr_data_18),
	.datac(\avl_rddata_local[13]~9_combout ),
	.datad(\csr_control_data[18]~q ),
	.cin(gnd),
	.combout(\rdata_comb[18]~139_combout ),
	.cout());
defparam \rdata_comb[18]~139 .lut_mask = 16'hE5E0;
defparam \rdata_comb[18]~139 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[18] (
	.clk(clk),
	.d(csr_wrdata[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[18]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[18] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[18] .power_up = "low";

dffeas \csr_wr_inst_data[18] (
	.clk(clk),
	.d(csr_wrdata[18]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(\csr_wr_inst_data[18]~q ),
	.prn(vcc));
defparam \csr_wr_inst_data[18] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[18] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[18]~140 (
	.dataa(avl_csr_address_3),
	.datab(\csr_flash_cmd_setting_data[18]~q ),
	.datac(avl_csr_address_0),
	.datad(\csr_wr_inst_data[18]~q ),
	.cin(gnd),
	.combout(\rdata_comb[18]~140_combout ),
	.cout());
defparam \rdata_comb[18]~140 .lut_mask = 16'hE5E0;
defparam \rdata_comb[18]~140 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[18]~141 (
	.dataa(csr_flash_cmd_wr_data_0_data_18),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[18]~140_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_18),
	.cin(gnd),
	.combout(\rdata_comb[18]~141_combout ),
	.cout());
defparam \rdata_comb[18]~141 .lut_mask = 16'hF838;
defparam \rdata_comb[18]~141 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[18]~142 (
	.dataa(\rdata_comb[18]~138_combout ),
	.datab(\avl_rddata_local[13]~8_combout ),
	.datac(\rdata_comb[18]~139_combout ),
	.datad(\rdata_comb[18]~141_combout ),
	.cin(gnd),
	.combout(\rdata_comb[18]~142_combout ),
	.cout());
defparam \rdata_comb[18]~142 .lut_mask = 16'hF838;
defparam \rdata_comb[18]~142 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[18]~143 (
	.dataa(\rdata_comb[18]~142_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avl_rddata_local[13]~10_combout ),
	.cin(gnd),
	.combout(\rdata_comb[18]~143_combout ),
	.cout());
defparam \rdata_comb[18]~143 .lut_mask = 16'h00AA;
defparam \rdata_comb[18]~143 .sum_lutc_input = "datac";

dffeas \csr_rd_inst_data[19] (
	.clk(clk),
	.d(csr_wrdata[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(\csr_rd_inst_data[19]~q ),
	.prn(vcc));
defparam \csr_rd_inst_data[19] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[19] .power_up = "low";

dffeas \csr_flash_cmd_rd_data_0_data[19] (
	.clk(clk),
	.d(out_rsp_data_19),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[19]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[19] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[19] .power_up = "low";

dffeas \csr_op_protocol_data[19] (
	.clk(clk),
	.d(csr_wrdata[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(\csr_op_protocol_data[19]~q ),
	.prn(vcc));
defparam \csr_op_protocol_data[19] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[19] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[19]~144 (
	.dataa(avl_csr_address_0),
	.datab(\csr_flash_cmd_rd_data_0_data[19]~q ),
	.datac(avl_csr_address_3),
	.datad(\csr_op_protocol_data[19]~q ),
	.cin(gnd),
	.combout(\rdata_comb[19]~144_combout ),
	.cout());
defparam \rdata_comb[19]~144 .lut_mask = 16'hE5E0;
defparam \rdata_comb[19]~144 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[19] (
	.clk(clk),
	.d(out_rsp_data_19),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[19]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[19] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[19] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[19]~145 (
	.dataa(\csr_rd_inst_data[19]~q ),
	.datab(avl_csr_address_0),
	.datac(\rdata_comb[19]~144_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[19]~q ),
	.cin(gnd),
	.combout(\rdata_comb[19]~145_combout ),
	.cout());
defparam \rdata_comb[19]~145 .lut_mask = 16'hF838;
defparam \rdata_comb[19]~145 .sum_lutc_input = "datac";

dffeas \csr_control_data[19] (
	.clk(clk),
	.d(csr_wrdata[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[19]~q ),
	.prn(vcc));
defparam \csr_control_data[19] .is_wysiwyg = "true";
defparam \csr_control_data[19] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[19]~146 (
	.dataa(\avl_rddata_local[13]~9_combout ),
	.datab(\rdata_comb[19]~145_combout ),
	.datac(\avl_rddata_local[13]~8_combout ),
	.datad(\csr_control_data[19]~q ),
	.cin(gnd),
	.combout(\rdata_comb[19]~146_combout ),
	.cout());
defparam \rdata_comb[19]~146 .lut_mask = 16'hE5E0;
defparam \rdata_comb[19]~146 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[19] (
	.clk(clk),
	.d(csr_wrdata[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[19]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[19] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[19] .power_up = "low";

dffeas \csr_wr_inst_data[19] (
	.clk(clk),
	.d(csr_wrdata[19]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(\csr_wr_inst_data[19]~q ),
	.prn(vcc));
defparam \csr_wr_inst_data[19] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[19] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[19]~147 (
	.dataa(avl_csr_address_3),
	.datab(\csr_flash_cmd_setting_data[19]~q ),
	.datac(avl_csr_address_0),
	.datad(\csr_wr_inst_data[19]~q ),
	.cin(gnd),
	.combout(\rdata_comb[19]~147_combout ),
	.cout());
defparam \rdata_comb[19]~147 .lut_mask = 16'hE5E0;
defparam \rdata_comb[19]~147 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[19]~148 (
	.dataa(csr_flash_cmd_wr_data_0_data_19),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[19]~147_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_19),
	.cin(gnd),
	.combout(\rdata_comb[19]~148_combout ),
	.cout());
defparam \rdata_comb[19]~148 .lut_mask = 16'hF838;
defparam \rdata_comb[19]~148 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[19]~149 (
	.dataa(csr_flash_cmd_addr_data_19),
	.datab(\avl_rddata_local[13]~9_combout ),
	.datac(\rdata_comb[19]~146_combout ),
	.datad(\rdata_comb[19]~148_combout ),
	.cin(gnd),
	.combout(\rdata_comb[19]~149_combout ),
	.cout());
defparam \rdata_comb[19]~149 .lut_mask = 16'hF838;
defparam \rdata_comb[19]~149 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[19]~150 (
	.dataa(\rdata_comb[19]~149_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avl_rddata_local[13]~10_combout ),
	.cin(gnd),
	.combout(\rdata_comb[19]~150_combout ),
	.cout());
defparam \rdata_comb[19]~150 .lut_mask = 16'h00AA;
defparam \rdata_comb[19]~150 .sum_lutc_input = "datac";

dffeas \csr_rd_inst_data[20] (
	.clk(clk),
	.d(csr_wrdata[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(\csr_rd_inst_data[20]~q ),
	.prn(vcc));
defparam \csr_rd_inst_data[20] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[20] .power_up = "low";

dffeas \csr_flash_cmd_rd_data_0_data[20] (
	.clk(clk),
	.d(out_rsp_data_20),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[20]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[20] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[20] .power_up = "low";

dffeas \csr_op_protocol_data[20] (
	.clk(clk),
	.d(csr_wrdata[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(\csr_op_protocol_data[20]~q ),
	.prn(vcc));
defparam \csr_op_protocol_data[20] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[20] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[20]~151 (
	.dataa(avl_csr_address_0),
	.datab(\csr_flash_cmd_rd_data_0_data[20]~q ),
	.datac(avl_csr_address_3),
	.datad(\csr_op_protocol_data[20]~q ),
	.cin(gnd),
	.combout(\rdata_comb[20]~151_combout ),
	.cout());
defparam \rdata_comb[20]~151 .lut_mask = 16'hE5E0;
defparam \rdata_comb[20]~151 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[20] (
	.clk(clk),
	.d(out_rsp_data_20),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[20]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[20] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[20] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[20]~152 (
	.dataa(\csr_rd_inst_data[20]~q ),
	.datab(avl_csr_address_0),
	.datac(\rdata_comb[20]~151_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[20]~q ),
	.cin(gnd),
	.combout(\rdata_comb[20]~152_combout ),
	.cout());
defparam \rdata_comb[20]~152 .lut_mask = 16'hF838;
defparam \rdata_comb[20]~152 .sum_lutc_input = "datac";

dffeas \csr_control_data[20] (
	.clk(clk),
	.d(csr_wrdata[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[20]~q ),
	.prn(vcc));
defparam \csr_control_data[20] .is_wysiwyg = "true";
defparam \csr_control_data[20] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[20]~153 (
	.dataa(\avl_rddata_local[13]~8_combout ),
	.datab(csr_flash_cmd_addr_data_20),
	.datac(\avl_rddata_local[13]~9_combout ),
	.datad(\csr_control_data[20]~q ),
	.cin(gnd),
	.combout(\rdata_comb[20]~153_combout ),
	.cout());
defparam \rdata_comb[20]~153 .lut_mask = 16'hE5E0;
defparam \rdata_comb[20]~153 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[20] (
	.clk(clk),
	.d(csr_wrdata[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[20]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[20] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[20] .power_up = "low";

dffeas \csr_wr_inst_data[20] (
	.clk(clk),
	.d(csr_wrdata[20]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(\csr_wr_inst_data[20]~q ),
	.prn(vcc));
defparam \csr_wr_inst_data[20] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[20] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[20]~154 (
	.dataa(avl_csr_address_3),
	.datab(\csr_flash_cmd_setting_data[20]~q ),
	.datac(avl_csr_address_0),
	.datad(\csr_wr_inst_data[20]~q ),
	.cin(gnd),
	.combout(\rdata_comb[20]~154_combout ),
	.cout());
defparam \rdata_comb[20]~154 .lut_mask = 16'hE5E0;
defparam \rdata_comb[20]~154 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[20]~155 (
	.dataa(csr_flash_cmd_wr_data_0_data_20),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[20]~154_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_20),
	.cin(gnd),
	.combout(\rdata_comb[20]~155_combout ),
	.cout());
defparam \rdata_comb[20]~155 .lut_mask = 16'hF838;
defparam \rdata_comb[20]~155 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[20]~156 (
	.dataa(\rdata_comb[20]~152_combout ),
	.datab(\avl_rddata_local[13]~8_combout ),
	.datac(\rdata_comb[20]~153_combout ),
	.datad(\rdata_comb[20]~155_combout ),
	.cin(gnd),
	.combout(\rdata_comb[20]~156_combout ),
	.cout());
defparam \rdata_comb[20]~156 .lut_mask = 16'hF838;
defparam \rdata_comb[20]~156 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[20]~157 (
	.dataa(\rdata_comb[20]~156_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avl_rddata_local[13]~10_combout ),
	.cin(gnd),
	.combout(\rdata_comb[20]~157_combout ),
	.cout());
defparam \rdata_comb[20]~157 .lut_mask = 16'h00AA;
defparam \rdata_comb[20]~157 .sum_lutc_input = "datac";

dffeas \csr_rd_inst_data[21] (
	.clk(clk),
	.d(csr_wrdata[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(\csr_rd_inst_data[21]~q ),
	.prn(vcc));
defparam \csr_rd_inst_data[21] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[21] .power_up = "low";

dffeas \csr_flash_cmd_rd_data_0_data[21] (
	.clk(clk),
	.d(out_rsp_data_21),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[21]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[21] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[21] .power_up = "low";

dffeas \csr_op_protocol_data[21] (
	.clk(clk),
	.d(csr_wrdata[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(\csr_op_protocol_data[21]~q ),
	.prn(vcc));
defparam \csr_op_protocol_data[21] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[21] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[21]~158 (
	.dataa(avl_csr_address_0),
	.datab(\csr_flash_cmd_rd_data_0_data[21]~q ),
	.datac(avl_csr_address_3),
	.datad(\csr_op_protocol_data[21]~q ),
	.cin(gnd),
	.combout(\rdata_comb[21]~158_combout ),
	.cout());
defparam \rdata_comb[21]~158 .lut_mask = 16'hE5E0;
defparam \rdata_comb[21]~158 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[21] (
	.clk(clk),
	.d(out_rsp_data_21),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[21]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[21] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[21] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[21]~159 (
	.dataa(\csr_rd_inst_data[21]~q ),
	.datab(avl_csr_address_0),
	.datac(\rdata_comb[21]~158_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[21]~q ),
	.cin(gnd),
	.combout(\rdata_comb[21]~159_combout ),
	.cout());
defparam \rdata_comb[21]~159 .lut_mask = 16'hF838;
defparam \rdata_comb[21]~159 .sum_lutc_input = "datac";

dffeas \csr_control_data[21] (
	.clk(clk),
	.d(csr_wrdata[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[21]~q ),
	.prn(vcc));
defparam \csr_control_data[21] .is_wysiwyg = "true";
defparam \csr_control_data[21] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[21]~160 (
	.dataa(\avl_rddata_local[13]~9_combout ),
	.datab(\rdata_comb[21]~159_combout ),
	.datac(\avl_rddata_local[13]~8_combout ),
	.datad(\csr_control_data[21]~q ),
	.cin(gnd),
	.combout(\rdata_comb[21]~160_combout ),
	.cout());
defparam \rdata_comb[21]~160 .lut_mask = 16'hE5E0;
defparam \rdata_comb[21]~160 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[21] (
	.clk(clk),
	.d(csr_wrdata[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[21]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[21] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[21] .power_up = "low";

dffeas \csr_wr_inst_data[21] (
	.clk(clk),
	.d(csr_wrdata[21]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(\csr_wr_inst_data[21]~q ),
	.prn(vcc));
defparam \csr_wr_inst_data[21] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[21] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[21]~161 (
	.dataa(avl_csr_address_3),
	.datab(\csr_flash_cmd_setting_data[21]~q ),
	.datac(avl_csr_address_0),
	.datad(\csr_wr_inst_data[21]~q ),
	.cin(gnd),
	.combout(\rdata_comb[21]~161_combout ),
	.cout());
defparam \rdata_comb[21]~161 .lut_mask = 16'hE5E0;
defparam \rdata_comb[21]~161 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[21]~162 (
	.dataa(csr_flash_cmd_wr_data_0_data_21),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[21]~161_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_21),
	.cin(gnd),
	.combout(\rdata_comb[21]~162_combout ),
	.cout());
defparam \rdata_comb[21]~162 .lut_mask = 16'hF838;
defparam \rdata_comb[21]~162 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[21]~163 (
	.dataa(csr_flash_cmd_addr_data_21),
	.datab(\avl_rddata_local[13]~9_combout ),
	.datac(\rdata_comb[21]~160_combout ),
	.datad(\rdata_comb[21]~162_combout ),
	.cin(gnd),
	.combout(\rdata_comb[21]~163_combout ),
	.cout());
defparam \rdata_comb[21]~163 .lut_mask = 16'hF838;
defparam \rdata_comb[21]~163 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[21]~164 (
	.dataa(\rdata_comb[21]~163_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avl_rddata_local[13]~10_combout ),
	.cin(gnd),
	.combout(\rdata_comb[21]~164_combout ),
	.cout());
defparam \rdata_comb[21]~164 .lut_mask = 16'h00AA;
defparam \rdata_comb[21]~164 .sum_lutc_input = "datac";

dffeas \csr_rd_inst_data[22] (
	.clk(clk),
	.d(csr_wrdata[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(\csr_rd_inst_data[22]~q ),
	.prn(vcc));
defparam \csr_rd_inst_data[22] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[22] .power_up = "low";

dffeas \csr_flash_cmd_rd_data_0_data[22] (
	.clk(clk),
	.d(out_rsp_data_22),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[22]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[22] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[22] .power_up = "low";

dffeas \csr_op_protocol_data[22] (
	.clk(clk),
	.d(csr_wrdata[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(\csr_op_protocol_data[22]~q ),
	.prn(vcc));
defparam \csr_op_protocol_data[22] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[22] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[22]~165 (
	.dataa(avl_csr_address_0),
	.datab(\csr_flash_cmd_rd_data_0_data[22]~q ),
	.datac(avl_csr_address_3),
	.datad(\csr_op_protocol_data[22]~q ),
	.cin(gnd),
	.combout(\rdata_comb[22]~165_combout ),
	.cout());
defparam \rdata_comb[22]~165 .lut_mask = 16'hE5E0;
defparam \rdata_comb[22]~165 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[22] (
	.clk(clk),
	.d(out_rsp_data_22),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[22]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[22] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[22] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[22]~166 (
	.dataa(\csr_rd_inst_data[22]~q ),
	.datab(avl_csr_address_0),
	.datac(\rdata_comb[22]~165_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[22]~q ),
	.cin(gnd),
	.combout(\rdata_comb[22]~166_combout ),
	.cout());
defparam \rdata_comb[22]~166 .lut_mask = 16'hF838;
defparam \rdata_comb[22]~166 .sum_lutc_input = "datac";

dffeas \csr_control_data[22] (
	.clk(clk),
	.d(csr_wrdata[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[22]~q ),
	.prn(vcc));
defparam \csr_control_data[22] .is_wysiwyg = "true";
defparam \csr_control_data[22] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[22]~167 (
	.dataa(\avl_rddata_local[13]~8_combout ),
	.datab(csr_flash_cmd_addr_data_22),
	.datac(\avl_rddata_local[13]~9_combout ),
	.datad(\csr_control_data[22]~q ),
	.cin(gnd),
	.combout(\rdata_comb[22]~167_combout ),
	.cout());
defparam \rdata_comb[22]~167 .lut_mask = 16'hE5E0;
defparam \rdata_comb[22]~167 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[22] (
	.clk(clk),
	.d(csr_wrdata[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[22]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[22] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[22] .power_up = "low";

dffeas \csr_wr_inst_data[22] (
	.clk(clk),
	.d(csr_wrdata[22]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(\csr_wr_inst_data[22]~q ),
	.prn(vcc));
defparam \csr_wr_inst_data[22] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[22] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[22]~168 (
	.dataa(avl_csr_address_3),
	.datab(\csr_flash_cmd_setting_data[22]~q ),
	.datac(avl_csr_address_0),
	.datad(\csr_wr_inst_data[22]~q ),
	.cin(gnd),
	.combout(\rdata_comb[22]~168_combout ),
	.cout());
defparam \rdata_comb[22]~168 .lut_mask = 16'hE5E0;
defparam \rdata_comb[22]~168 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[22]~169 (
	.dataa(csr_flash_cmd_wr_data_0_data_22),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[22]~168_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_22),
	.cin(gnd),
	.combout(\rdata_comb[22]~169_combout ),
	.cout());
defparam \rdata_comb[22]~169 .lut_mask = 16'hF838;
defparam \rdata_comb[22]~169 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[22]~170 (
	.dataa(\rdata_comb[22]~166_combout ),
	.datab(\avl_rddata_local[13]~8_combout ),
	.datac(\rdata_comb[22]~167_combout ),
	.datad(\rdata_comb[22]~169_combout ),
	.cin(gnd),
	.combout(\rdata_comb[22]~170_combout ),
	.cout());
defparam \rdata_comb[22]~170 .lut_mask = 16'hF838;
defparam \rdata_comb[22]~170 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[22]~171 (
	.dataa(\rdata_comb[22]~170_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avl_rddata_local[13]~10_combout ),
	.cin(gnd),
	.combout(\rdata_comb[22]~171_combout ),
	.cout());
defparam \rdata_comb[22]~171 .lut_mask = 16'h00AA;
defparam \rdata_comb[22]~171 .sum_lutc_input = "datac";

dffeas \csr_rd_inst_data[23] (
	.clk(clk),
	.d(csr_wrdata[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(\csr_rd_inst_data[23]~q ),
	.prn(vcc));
defparam \csr_rd_inst_data[23] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[23] .power_up = "low";

dffeas \csr_flash_cmd_rd_data_0_data[23] (
	.clk(clk),
	.d(out_rsp_data_23),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[23]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[23] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[23] .power_up = "low";

dffeas \csr_op_protocol_data[23] (
	.clk(clk),
	.d(csr_wrdata[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(\csr_op_protocol_data[23]~q ),
	.prn(vcc));
defparam \csr_op_protocol_data[23] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[23] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[23]~172 (
	.dataa(avl_csr_address_0),
	.datab(\csr_flash_cmd_rd_data_0_data[23]~q ),
	.datac(avl_csr_address_3),
	.datad(\csr_op_protocol_data[23]~q ),
	.cin(gnd),
	.combout(\rdata_comb[23]~172_combout ),
	.cout());
defparam \rdata_comb[23]~172 .lut_mask = 16'hE5E0;
defparam \rdata_comb[23]~172 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[23] (
	.clk(clk),
	.d(out_rsp_data_23),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[23]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[23] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[23] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[23]~173 (
	.dataa(\csr_rd_inst_data[23]~q ),
	.datab(avl_csr_address_0),
	.datac(\rdata_comb[23]~172_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[23]~q ),
	.cin(gnd),
	.combout(\rdata_comb[23]~173_combout ),
	.cout());
defparam \rdata_comb[23]~173 .lut_mask = 16'hF838;
defparam \rdata_comb[23]~173 .sum_lutc_input = "datac";

dffeas \csr_control_data[23] (
	.clk(clk),
	.d(csr_wrdata[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[23]~q ),
	.prn(vcc));
defparam \csr_control_data[23] .is_wysiwyg = "true";
defparam \csr_control_data[23] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[23]~174 (
	.dataa(\avl_rddata_local[13]~9_combout ),
	.datab(\rdata_comb[23]~173_combout ),
	.datac(\avl_rddata_local[13]~8_combout ),
	.datad(\csr_control_data[23]~q ),
	.cin(gnd),
	.combout(\rdata_comb[23]~174_combout ),
	.cout());
defparam \rdata_comb[23]~174 .lut_mask = 16'hE5E0;
defparam \rdata_comb[23]~174 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[23] (
	.clk(clk),
	.d(csr_wrdata[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[23]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[23] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[23] .power_up = "low";

dffeas \csr_wr_inst_data[23] (
	.clk(clk),
	.d(csr_wrdata[23]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(\csr_wr_inst_data[23]~q ),
	.prn(vcc));
defparam \csr_wr_inst_data[23] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[23] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[23]~175 (
	.dataa(avl_csr_address_3),
	.datab(\csr_flash_cmd_setting_data[23]~q ),
	.datac(avl_csr_address_0),
	.datad(\csr_wr_inst_data[23]~q ),
	.cin(gnd),
	.combout(\rdata_comb[23]~175_combout ),
	.cout());
defparam \rdata_comb[23]~175 .lut_mask = 16'hE5E0;
defparam \rdata_comb[23]~175 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[23]~176 (
	.dataa(csr_flash_cmd_wr_data_0_data_23),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[23]~175_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_23),
	.cin(gnd),
	.combout(\rdata_comb[23]~176_combout ),
	.cout());
defparam \rdata_comb[23]~176 .lut_mask = 16'hF838;
defparam \rdata_comb[23]~176 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[23]~177 (
	.dataa(csr_flash_cmd_addr_data_23),
	.datab(\avl_rddata_local[13]~9_combout ),
	.datac(\rdata_comb[23]~174_combout ),
	.datad(\rdata_comb[23]~176_combout ),
	.cin(gnd),
	.combout(\rdata_comb[23]~177_combout ),
	.cout());
defparam \rdata_comb[23]~177 .lut_mask = 16'hF838;
defparam \rdata_comb[23]~177 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[23]~178 (
	.dataa(\rdata_comb[23]~177_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avl_rddata_local[13]~10_combout ),
	.cin(gnd),
	.combout(\rdata_comb[23]~178_combout ),
	.cout());
defparam \rdata_comb[23]~178 .lut_mask = 16'h00AA;
defparam \rdata_comb[23]~178 .sum_lutc_input = "datac";

dffeas \csr_rd_inst_data[24] (
	.clk(clk),
	.d(csr_wrdata[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(\csr_rd_inst_data[24]~q ),
	.prn(vcc));
defparam \csr_rd_inst_data[24] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[24] .power_up = "low";

dffeas \csr_flash_cmd_rd_data_0_data[24] (
	.clk(clk),
	.d(out_rsp_data_24),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[24]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[24] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[24] .power_up = "low";

dffeas \csr_op_protocol_data[24] (
	.clk(clk),
	.d(csr_wrdata[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(\csr_op_protocol_data[24]~q ),
	.prn(vcc));
defparam \csr_op_protocol_data[24] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[24] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[24]~179 (
	.dataa(avl_csr_address_0),
	.datab(\csr_flash_cmd_rd_data_0_data[24]~q ),
	.datac(avl_csr_address_3),
	.datad(\csr_op_protocol_data[24]~q ),
	.cin(gnd),
	.combout(\rdata_comb[24]~179_combout ),
	.cout());
defparam \rdata_comb[24]~179 .lut_mask = 16'hE5E0;
defparam \rdata_comb[24]~179 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[24] (
	.clk(clk),
	.d(out_rsp_data_24),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[24]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[24] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[24] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[24]~180 (
	.dataa(\csr_rd_inst_data[24]~q ),
	.datab(avl_csr_address_0),
	.datac(\rdata_comb[24]~179_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[24]~q ),
	.cin(gnd),
	.combout(\rdata_comb[24]~180_combout ),
	.cout());
defparam \rdata_comb[24]~180 .lut_mask = 16'hF838;
defparam \rdata_comb[24]~180 .sum_lutc_input = "datac";

dffeas \csr_control_data[24] (
	.clk(clk),
	.d(csr_wrdata[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[24]~q ),
	.prn(vcc));
defparam \csr_control_data[24] .is_wysiwyg = "true";
defparam \csr_control_data[24] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[24]~181 (
	.dataa(\avl_rddata_local[13]~8_combout ),
	.datab(csr_flash_cmd_addr_data_24),
	.datac(\avl_rddata_local[13]~9_combout ),
	.datad(\csr_control_data[24]~q ),
	.cin(gnd),
	.combout(\rdata_comb[24]~181_combout ),
	.cout());
defparam \rdata_comb[24]~181 .lut_mask = 16'hE5E0;
defparam \rdata_comb[24]~181 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[24] (
	.clk(clk),
	.d(csr_wrdata[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[24]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[24] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[24] .power_up = "low";

dffeas \csr_wr_inst_data[24] (
	.clk(clk),
	.d(csr_wrdata[24]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(\csr_wr_inst_data[24]~q ),
	.prn(vcc));
defparam \csr_wr_inst_data[24] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[24] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[24]~182 (
	.dataa(avl_csr_address_3),
	.datab(\csr_flash_cmd_setting_data[24]~q ),
	.datac(avl_csr_address_0),
	.datad(\csr_wr_inst_data[24]~q ),
	.cin(gnd),
	.combout(\rdata_comb[24]~182_combout ),
	.cout());
defparam \rdata_comb[24]~182 .lut_mask = 16'hE5E0;
defparam \rdata_comb[24]~182 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[24]~183 (
	.dataa(csr_flash_cmd_wr_data_0_data_24),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[24]~182_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_24),
	.cin(gnd),
	.combout(\rdata_comb[24]~183_combout ),
	.cout());
defparam \rdata_comb[24]~183 .lut_mask = 16'hF838;
defparam \rdata_comb[24]~183 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[24]~184 (
	.dataa(\rdata_comb[24]~180_combout ),
	.datab(\avl_rddata_local[13]~8_combout ),
	.datac(\rdata_comb[24]~181_combout ),
	.datad(\rdata_comb[24]~183_combout ),
	.cin(gnd),
	.combout(\rdata_comb[24]~184_combout ),
	.cout());
defparam \rdata_comb[24]~184 .lut_mask = 16'hF838;
defparam \rdata_comb[24]~184 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[24]~185 (
	.dataa(\rdata_comb[24]~184_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avl_rddata_local[13]~10_combout ),
	.cin(gnd),
	.combout(\rdata_comb[24]~185_combout ),
	.cout());
defparam \rdata_comb[24]~185 .lut_mask = 16'h00AA;
defparam \rdata_comb[24]~185 .sum_lutc_input = "datac";

dffeas \csr_rd_inst_data[25] (
	.clk(clk),
	.d(csr_wrdata[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(\csr_rd_inst_data[25]~q ),
	.prn(vcc));
defparam \csr_rd_inst_data[25] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[25] .power_up = "low";

dffeas \csr_flash_cmd_rd_data_0_data[25] (
	.clk(clk),
	.d(out_rsp_data_25),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[25]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[25] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[25] .power_up = "low";

dffeas \csr_op_protocol_data[25] (
	.clk(clk),
	.d(csr_wrdata[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(\csr_op_protocol_data[25]~q ),
	.prn(vcc));
defparam \csr_op_protocol_data[25] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[25] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[25]~186 (
	.dataa(avl_csr_address_0),
	.datab(\csr_flash_cmd_rd_data_0_data[25]~q ),
	.datac(avl_csr_address_3),
	.datad(\csr_op_protocol_data[25]~q ),
	.cin(gnd),
	.combout(\rdata_comb[25]~186_combout ),
	.cout());
defparam \rdata_comb[25]~186 .lut_mask = 16'hE5E0;
defparam \rdata_comb[25]~186 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[25] (
	.clk(clk),
	.d(out_rsp_data_25),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[25]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[25] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[25] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[25]~187 (
	.dataa(\csr_rd_inst_data[25]~q ),
	.datab(avl_csr_address_0),
	.datac(\rdata_comb[25]~186_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[25]~q ),
	.cin(gnd),
	.combout(\rdata_comb[25]~187_combout ),
	.cout());
defparam \rdata_comb[25]~187 .lut_mask = 16'hF838;
defparam \rdata_comb[25]~187 .sum_lutc_input = "datac";

dffeas \csr_control_data[25] (
	.clk(clk),
	.d(csr_wrdata[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[25]~q ),
	.prn(vcc));
defparam \csr_control_data[25] .is_wysiwyg = "true";
defparam \csr_control_data[25] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[25]~188 (
	.dataa(\avl_rddata_local[13]~9_combout ),
	.datab(\rdata_comb[25]~187_combout ),
	.datac(\avl_rddata_local[13]~8_combout ),
	.datad(\csr_control_data[25]~q ),
	.cin(gnd),
	.combout(\rdata_comb[25]~188_combout ),
	.cout());
defparam \rdata_comb[25]~188 .lut_mask = 16'hE5E0;
defparam \rdata_comb[25]~188 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[25] (
	.clk(clk),
	.d(csr_wrdata[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[25]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[25] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[25] .power_up = "low";

dffeas \csr_wr_inst_data[25] (
	.clk(clk),
	.d(csr_wrdata[25]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(\csr_wr_inst_data[25]~q ),
	.prn(vcc));
defparam \csr_wr_inst_data[25] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[25] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[25]~189 (
	.dataa(avl_csr_address_3),
	.datab(\csr_flash_cmd_setting_data[25]~q ),
	.datac(avl_csr_address_0),
	.datad(\csr_wr_inst_data[25]~q ),
	.cin(gnd),
	.combout(\rdata_comb[25]~189_combout ),
	.cout());
defparam \rdata_comb[25]~189 .lut_mask = 16'hE5E0;
defparam \rdata_comb[25]~189 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[25]~190 (
	.dataa(csr_flash_cmd_wr_data_0_data_25),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[25]~189_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_25),
	.cin(gnd),
	.combout(\rdata_comb[25]~190_combout ),
	.cout());
defparam \rdata_comb[25]~190 .lut_mask = 16'hF838;
defparam \rdata_comb[25]~190 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[25]~191 (
	.dataa(csr_flash_cmd_addr_data_25),
	.datab(\avl_rddata_local[13]~9_combout ),
	.datac(\rdata_comb[25]~188_combout ),
	.datad(\rdata_comb[25]~190_combout ),
	.cin(gnd),
	.combout(\rdata_comb[25]~191_combout ),
	.cout());
defparam \rdata_comb[25]~191 .lut_mask = 16'hF838;
defparam \rdata_comb[25]~191 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[25]~192 (
	.dataa(\rdata_comb[25]~191_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avl_rddata_local[13]~10_combout ),
	.cin(gnd),
	.combout(\rdata_comb[25]~192_combout ),
	.cout());
defparam \rdata_comb[25]~192 .lut_mask = 16'h00AA;
defparam \rdata_comb[25]~192 .sum_lutc_input = "datac";

dffeas \csr_rd_inst_data[26] (
	.clk(clk),
	.d(csr_wrdata[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(\csr_rd_inst_data[26]~q ),
	.prn(vcc));
defparam \csr_rd_inst_data[26] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[26] .power_up = "low";

dffeas \csr_flash_cmd_rd_data_0_data[26] (
	.clk(clk),
	.d(out_rsp_data_26),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[26]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[26] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[26] .power_up = "low";

dffeas \csr_op_protocol_data[26] (
	.clk(clk),
	.d(csr_wrdata[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(\csr_op_protocol_data[26]~q ),
	.prn(vcc));
defparam \csr_op_protocol_data[26] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[26] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[26]~193 (
	.dataa(avl_csr_address_0),
	.datab(\csr_flash_cmd_rd_data_0_data[26]~q ),
	.datac(avl_csr_address_3),
	.datad(\csr_op_protocol_data[26]~q ),
	.cin(gnd),
	.combout(\rdata_comb[26]~193_combout ),
	.cout());
defparam \rdata_comb[26]~193 .lut_mask = 16'hE5E0;
defparam \rdata_comb[26]~193 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[26] (
	.clk(clk),
	.d(out_rsp_data_26),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[26]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[26] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[26] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[26]~194 (
	.dataa(\csr_rd_inst_data[26]~q ),
	.datab(avl_csr_address_0),
	.datac(\rdata_comb[26]~193_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[26]~q ),
	.cin(gnd),
	.combout(\rdata_comb[26]~194_combout ),
	.cout());
defparam \rdata_comb[26]~194 .lut_mask = 16'hF838;
defparam \rdata_comb[26]~194 .sum_lutc_input = "datac";

dffeas \csr_control_data[26] (
	.clk(clk),
	.d(csr_wrdata[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[26]~q ),
	.prn(vcc));
defparam \csr_control_data[26] .is_wysiwyg = "true";
defparam \csr_control_data[26] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[26]~195 (
	.dataa(\avl_rddata_local[13]~8_combout ),
	.datab(csr_flash_cmd_addr_data_26),
	.datac(\avl_rddata_local[13]~9_combout ),
	.datad(\csr_control_data[26]~q ),
	.cin(gnd),
	.combout(\rdata_comb[26]~195_combout ),
	.cout());
defparam \rdata_comb[26]~195 .lut_mask = 16'hE5E0;
defparam \rdata_comb[26]~195 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[26] (
	.clk(clk),
	.d(csr_wrdata[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[26]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[26] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[26] .power_up = "low";

dffeas \csr_wr_inst_data[26] (
	.clk(clk),
	.d(csr_wrdata[26]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(\csr_wr_inst_data[26]~q ),
	.prn(vcc));
defparam \csr_wr_inst_data[26] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[26] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[26]~196 (
	.dataa(avl_csr_address_3),
	.datab(\csr_flash_cmd_setting_data[26]~q ),
	.datac(avl_csr_address_0),
	.datad(\csr_wr_inst_data[26]~q ),
	.cin(gnd),
	.combout(\rdata_comb[26]~196_combout ),
	.cout());
defparam \rdata_comb[26]~196 .lut_mask = 16'hE5E0;
defparam \rdata_comb[26]~196 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[26]~197 (
	.dataa(csr_flash_cmd_wr_data_0_data_26),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[26]~196_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_26),
	.cin(gnd),
	.combout(\rdata_comb[26]~197_combout ),
	.cout());
defparam \rdata_comb[26]~197 .lut_mask = 16'hF838;
defparam \rdata_comb[26]~197 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[26]~198 (
	.dataa(\rdata_comb[26]~194_combout ),
	.datab(\avl_rddata_local[13]~8_combout ),
	.datac(\rdata_comb[26]~195_combout ),
	.datad(\rdata_comb[26]~197_combout ),
	.cin(gnd),
	.combout(\rdata_comb[26]~198_combout ),
	.cout());
defparam \rdata_comb[26]~198 .lut_mask = 16'hF838;
defparam \rdata_comb[26]~198 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[26]~199 (
	.dataa(\rdata_comb[26]~198_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avl_rddata_local[13]~10_combout ),
	.cin(gnd),
	.combout(\rdata_comb[26]~199_combout ),
	.cout());
defparam \rdata_comb[26]~199 .lut_mask = 16'h00AA;
defparam \rdata_comb[26]~199 .sum_lutc_input = "datac";

dffeas \csr_rd_inst_data[27] (
	.clk(clk),
	.d(csr_wrdata[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(\csr_rd_inst_data[27]~q ),
	.prn(vcc));
defparam \csr_rd_inst_data[27] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[27] .power_up = "low";

dffeas \csr_flash_cmd_rd_data_0_data[27] (
	.clk(clk),
	.d(out_rsp_data_27),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[27]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[27] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[27] .power_up = "low";

dffeas \csr_op_protocol_data[27] (
	.clk(clk),
	.d(csr_wrdata[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(\csr_op_protocol_data[27]~q ),
	.prn(vcc));
defparam \csr_op_protocol_data[27] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[27] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[27]~200 (
	.dataa(avl_csr_address_0),
	.datab(\csr_flash_cmd_rd_data_0_data[27]~q ),
	.datac(avl_csr_address_3),
	.datad(\csr_op_protocol_data[27]~q ),
	.cin(gnd),
	.combout(\rdata_comb[27]~200_combout ),
	.cout());
defparam \rdata_comb[27]~200 .lut_mask = 16'hE5E0;
defparam \rdata_comb[27]~200 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[27] (
	.clk(clk),
	.d(out_rsp_data_27),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[27]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[27] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[27] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[27]~201 (
	.dataa(\csr_rd_inst_data[27]~q ),
	.datab(avl_csr_address_0),
	.datac(\rdata_comb[27]~200_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[27]~q ),
	.cin(gnd),
	.combout(\rdata_comb[27]~201_combout ),
	.cout());
defparam \rdata_comb[27]~201 .lut_mask = 16'hF838;
defparam \rdata_comb[27]~201 .sum_lutc_input = "datac";

dffeas \csr_control_data[27] (
	.clk(clk),
	.d(csr_wrdata[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[27]~q ),
	.prn(vcc));
defparam \csr_control_data[27] .is_wysiwyg = "true";
defparam \csr_control_data[27] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[27]~202 (
	.dataa(\avl_rddata_local[13]~9_combout ),
	.datab(\rdata_comb[27]~201_combout ),
	.datac(\avl_rddata_local[13]~8_combout ),
	.datad(\csr_control_data[27]~q ),
	.cin(gnd),
	.combout(\rdata_comb[27]~202_combout ),
	.cout());
defparam \rdata_comb[27]~202 .lut_mask = 16'hE5E0;
defparam \rdata_comb[27]~202 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[27] (
	.clk(clk),
	.d(csr_wrdata[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[27]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[27] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[27] .power_up = "low";

dffeas \csr_wr_inst_data[27] (
	.clk(clk),
	.d(csr_wrdata[27]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(\csr_wr_inst_data[27]~q ),
	.prn(vcc));
defparam \csr_wr_inst_data[27] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[27] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[27]~203 (
	.dataa(avl_csr_address_3),
	.datab(\csr_flash_cmd_setting_data[27]~q ),
	.datac(avl_csr_address_0),
	.datad(\csr_wr_inst_data[27]~q ),
	.cin(gnd),
	.combout(\rdata_comb[27]~203_combout ),
	.cout());
defparam \rdata_comb[27]~203 .lut_mask = 16'hE5E0;
defparam \rdata_comb[27]~203 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[27]~204 (
	.dataa(csr_flash_cmd_wr_data_0_data_27),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[27]~203_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_27),
	.cin(gnd),
	.combout(\rdata_comb[27]~204_combout ),
	.cout());
defparam \rdata_comb[27]~204 .lut_mask = 16'hF838;
defparam \rdata_comb[27]~204 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[27]~205 (
	.dataa(csr_flash_cmd_addr_data_27),
	.datab(\avl_rddata_local[13]~9_combout ),
	.datac(\rdata_comb[27]~202_combout ),
	.datad(\rdata_comb[27]~204_combout ),
	.cin(gnd),
	.combout(\rdata_comb[27]~205_combout ),
	.cout());
defparam \rdata_comb[27]~205 .lut_mask = 16'hF838;
defparam \rdata_comb[27]~205 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[27]~206 (
	.dataa(\rdata_comb[27]~205_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avl_rddata_local[13]~10_combout ),
	.cin(gnd),
	.combout(\rdata_comb[27]~206_combout ),
	.cout());
defparam \rdata_comb[27]~206 .lut_mask = 16'h00AA;
defparam \rdata_comb[27]~206 .sum_lutc_input = "datac";

dffeas \csr_rd_inst_data[28] (
	.clk(clk),
	.d(csr_wrdata[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(\csr_rd_inst_data[28]~q ),
	.prn(vcc));
defparam \csr_rd_inst_data[28] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[28] .power_up = "low";

dffeas \csr_flash_cmd_rd_data_0_data[28] (
	.clk(clk),
	.d(out_rsp_data_28),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[28]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[28] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[28] .power_up = "low";

dffeas \csr_op_protocol_data[28] (
	.clk(clk),
	.d(csr_wrdata[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(\csr_op_protocol_data[28]~q ),
	.prn(vcc));
defparam \csr_op_protocol_data[28] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[28] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[28]~207 (
	.dataa(avl_csr_address_0),
	.datab(\csr_flash_cmd_rd_data_0_data[28]~q ),
	.datac(avl_csr_address_3),
	.datad(\csr_op_protocol_data[28]~q ),
	.cin(gnd),
	.combout(\rdata_comb[28]~207_combout ),
	.cout());
defparam \rdata_comb[28]~207 .lut_mask = 16'hE5E0;
defparam \rdata_comb[28]~207 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[28] (
	.clk(clk),
	.d(out_rsp_data_28),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[28]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[28] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[28] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[28]~208 (
	.dataa(\csr_rd_inst_data[28]~q ),
	.datab(avl_csr_address_0),
	.datac(\rdata_comb[28]~207_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[28]~q ),
	.cin(gnd),
	.combout(\rdata_comb[28]~208_combout ),
	.cout());
defparam \rdata_comb[28]~208 .lut_mask = 16'hF838;
defparam \rdata_comb[28]~208 .sum_lutc_input = "datac";

dffeas \csr_control_data[28] (
	.clk(clk),
	.d(csr_wrdata[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[28]~q ),
	.prn(vcc));
defparam \csr_control_data[28] .is_wysiwyg = "true";
defparam \csr_control_data[28] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[28]~209 (
	.dataa(\avl_rddata_local[13]~8_combout ),
	.datab(csr_flash_cmd_addr_data_28),
	.datac(\avl_rddata_local[13]~9_combout ),
	.datad(\csr_control_data[28]~q ),
	.cin(gnd),
	.combout(\rdata_comb[28]~209_combout ),
	.cout());
defparam \rdata_comb[28]~209 .lut_mask = 16'hE5E0;
defparam \rdata_comb[28]~209 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[28] (
	.clk(clk),
	.d(csr_wrdata[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[28]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[28] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[28] .power_up = "low";

dffeas \csr_wr_inst_data[28] (
	.clk(clk),
	.d(csr_wrdata[28]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(\csr_wr_inst_data[28]~q ),
	.prn(vcc));
defparam \csr_wr_inst_data[28] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[28] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[28]~210 (
	.dataa(avl_csr_address_3),
	.datab(\csr_flash_cmd_setting_data[28]~q ),
	.datac(avl_csr_address_0),
	.datad(\csr_wr_inst_data[28]~q ),
	.cin(gnd),
	.combout(\rdata_comb[28]~210_combout ),
	.cout());
defparam \rdata_comb[28]~210 .lut_mask = 16'hE5E0;
defparam \rdata_comb[28]~210 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[28]~211 (
	.dataa(csr_flash_cmd_wr_data_0_data_28),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[28]~210_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_28),
	.cin(gnd),
	.combout(\rdata_comb[28]~211_combout ),
	.cout());
defparam \rdata_comb[28]~211 .lut_mask = 16'hF838;
defparam \rdata_comb[28]~211 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[28]~212 (
	.dataa(\rdata_comb[28]~208_combout ),
	.datab(\avl_rddata_local[13]~8_combout ),
	.datac(\rdata_comb[28]~209_combout ),
	.datad(\rdata_comb[28]~211_combout ),
	.cin(gnd),
	.combout(\rdata_comb[28]~212_combout ),
	.cout());
defparam \rdata_comb[28]~212 .lut_mask = 16'hF838;
defparam \rdata_comb[28]~212 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[28]~213 (
	.dataa(\rdata_comb[28]~212_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avl_rddata_local[13]~10_combout ),
	.cin(gnd),
	.combout(\rdata_comb[28]~213_combout ),
	.cout());
defparam \rdata_comb[28]~213 .lut_mask = 16'h00AA;
defparam \rdata_comb[28]~213 .sum_lutc_input = "datac";

dffeas \csr_rd_inst_data[29] (
	.clk(clk),
	.d(csr_wrdata[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(\csr_rd_inst_data[29]~q ),
	.prn(vcc));
defparam \csr_rd_inst_data[29] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[29] .power_up = "low";

dffeas \csr_flash_cmd_rd_data_0_data[29] (
	.clk(clk),
	.d(out_rsp_data_29),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[29]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[29] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[29] .power_up = "low";

dffeas \csr_op_protocol_data[29] (
	.clk(clk),
	.d(csr_wrdata[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(\csr_op_protocol_data[29]~q ),
	.prn(vcc));
defparam \csr_op_protocol_data[29] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[29] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[29]~214 (
	.dataa(avl_csr_address_0),
	.datab(\csr_flash_cmd_rd_data_0_data[29]~q ),
	.datac(avl_csr_address_3),
	.datad(\csr_op_protocol_data[29]~q ),
	.cin(gnd),
	.combout(\rdata_comb[29]~214_combout ),
	.cout());
defparam \rdata_comb[29]~214 .lut_mask = 16'hE5E0;
defparam \rdata_comb[29]~214 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[29] (
	.clk(clk),
	.d(out_rsp_data_29),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[29]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[29] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[29] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[29]~215 (
	.dataa(\csr_rd_inst_data[29]~q ),
	.datab(avl_csr_address_0),
	.datac(\rdata_comb[29]~214_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[29]~q ),
	.cin(gnd),
	.combout(\rdata_comb[29]~215_combout ),
	.cout());
defparam \rdata_comb[29]~215 .lut_mask = 16'hF838;
defparam \rdata_comb[29]~215 .sum_lutc_input = "datac";

dffeas \csr_control_data[29] (
	.clk(clk),
	.d(csr_wrdata[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[29]~q ),
	.prn(vcc));
defparam \csr_control_data[29] .is_wysiwyg = "true";
defparam \csr_control_data[29] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[29]~216 (
	.dataa(\avl_rddata_local[13]~9_combout ),
	.datab(\rdata_comb[29]~215_combout ),
	.datac(\avl_rddata_local[13]~8_combout ),
	.datad(\csr_control_data[29]~q ),
	.cin(gnd),
	.combout(\rdata_comb[29]~216_combout ),
	.cout());
defparam \rdata_comb[29]~216 .lut_mask = 16'hE5E0;
defparam \rdata_comb[29]~216 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[29] (
	.clk(clk),
	.d(csr_wrdata[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[29]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[29] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[29] .power_up = "low";

dffeas \csr_wr_inst_data[29] (
	.clk(clk),
	.d(csr_wrdata[29]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(\csr_wr_inst_data[29]~q ),
	.prn(vcc));
defparam \csr_wr_inst_data[29] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[29] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[29]~217 (
	.dataa(avl_csr_address_3),
	.datab(\csr_flash_cmd_setting_data[29]~q ),
	.datac(avl_csr_address_0),
	.datad(\csr_wr_inst_data[29]~q ),
	.cin(gnd),
	.combout(\rdata_comb[29]~217_combout ),
	.cout());
defparam \rdata_comb[29]~217 .lut_mask = 16'hE5E0;
defparam \rdata_comb[29]~217 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[29]~218 (
	.dataa(csr_flash_cmd_wr_data_0_data_29),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[29]~217_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_29),
	.cin(gnd),
	.combout(\rdata_comb[29]~218_combout ),
	.cout());
defparam \rdata_comb[29]~218 .lut_mask = 16'hF838;
defparam \rdata_comb[29]~218 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[29]~219 (
	.dataa(csr_flash_cmd_addr_data_29),
	.datab(\avl_rddata_local[13]~9_combout ),
	.datac(\rdata_comb[29]~216_combout ),
	.datad(\rdata_comb[29]~218_combout ),
	.cin(gnd),
	.combout(\rdata_comb[29]~219_combout ),
	.cout());
defparam \rdata_comb[29]~219 .lut_mask = 16'hF838;
defparam \rdata_comb[29]~219 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[29]~220 (
	.dataa(\rdata_comb[29]~219_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avl_rddata_local[13]~10_combout ),
	.cin(gnd),
	.combout(\rdata_comb[29]~220_combout ),
	.cout());
defparam \rdata_comb[29]~220 .lut_mask = 16'h00AA;
defparam \rdata_comb[29]~220 .sum_lutc_input = "datac";

dffeas \csr_rd_inst_data[30] (
	.clk(clk),
	.d(csr_wrdata[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(\csr_rd_inst_data[30]~q ),
	.prn(vcc));
defparam \csr_rd_inst_data[30] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[30] .power_up = "low";

dffeas \csr_flash_cmd_rd_data_0_data[30] (
	.clk(clk),
	.d(out_rsp_data_30),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[30]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[30] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[30] .power_up = "low";

dffeas \csr_op_protocol_data[30] (
	.clk(clk),
	.d(csr_wrdata[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(\csr_op_protocol_data[30]~q ),
	.prn(vcc));
defparam \csr_op_protocol_data[30] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[30] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[30]~221 (
	.dataa(avl_csr_address_0),
	.datab(\csr_flash_cmd_rd_data_0_data[30]~q ),
	.datac(avl_csr_address_3),
	.datad(\csr_op_protocol_data[30]~q ),
	.cin(gnd),
	.combout(\rdata_comb[30]~221_combout ),
	.cout());
defparam \rdata_comb[30]~221 .lut_mask = 16'hE5E0;
defparam \rdata_comb[30]~221 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[30] (
	.clk(clk),
	.d(out_rsp_data_30),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[30]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[30] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[30] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[30]~222 (
	.dataa(\csr_rd_inst_data[30]~q ),
	.datab(avl_csr_address_0),
	.datac(\rdata_comb[30]~221_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[30]~q ),
	.cin(gnd),
	.combout(\rdata_comb[30]~222_combout ),
	.cout());
defparam \rdata_comb[30]~222 .lut_mask = 16'hF838;
defparam \rdata_comb[30]~222 .sum_lutc_input = "datac";

dffeas \csr_control_data[30] (
	.clk(clk),
	.d(csr_wrdata[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[30]~q ),
	.prn(vcc));
defparam \csr_control_data[30] .is_wysiwyg = "true";
defparam \csr_control_data[30] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[30]~223 (
	.dataa(\avl_rddata_local[13]~8_combout ),
	.datab(csr_flash_cmd_addr_data_30),
	.datac(\avl_rddata_local[13]~9_combout ),
	.datad(\csr_control_data[30]~q ),
	.cin(gnd),
	.combout(\rdata_comb[30]~223_combout ),
	.cout());
defparam \rdata_comb[30]~223 .lut_mask = 16'hE5E0;
defparam \rdata_comb[30]~223 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[30] (
	.clk(clk),
	.d(csr_wrdata[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[30]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[30] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[30] .power_up = "low";

dffeas \csr_wr_inst_data[30] (
	.clk(clk),
	.d(csr_wrdata[30]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(\csr_wr_inst_data[30]~q ),
	.prn(vcc));
defparam \csr_wr_inst_data[30] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[30] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[30]~224 (
	.dataa(avl_csr_address_3),
	.datab(\csr_flash_cmd_setting_data[30]~q ),
	.datac(avl_csr_address_0),
	.datad(\csr_wr_inst_data[30]~q ),
	.cin(gnd),
	.combout(\rdata_comb[30]~224_combout ),
	.cout());
defparam \rdata_comb[30]~224 .lut_mask = 16'hE5E0;
defparam \rdata_comb[30]~224 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[30]~225 (
	.dataa(csr_flash_cmd_wr_data_0_data_30),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[30]~224_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_30),
	.cin(gnd),
	.combout(\rdata_comb[30]~225_combout ),
	.cout());
defparam \rdata_comb[30]~225 .lut_mask = 16'hF838;
defparam \rdata_comb[30]~225 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[30]~226 (
	.dataa(\rdata_comb[30]~222_combout ),
	.datab(\avl_rddata_local[13]~8_combout ),
	.datac(\rdata_comb[30]~223_combout ),
	.datad(\rdata_comb[30]~225_combout ),
	.cin(gnd),
	.combout(\rdata_comb[30]~226_combout ),
	.cout());
defparam \rdata_comb[30]~226 .lut_mask = 16'hF838;
defparam \rdata_comb[30]~226 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[30]~227 (
	.dataa(\rdata_comb[30]~226_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avl_rddata_local[13]~10_combout ),
	.cin(gnd),
	.combout(\rdata_comb[30]~227_combout ),
	.cout());
defparam \rdata_comb[30]~227 .lut_mask = 16'h00AA;
defparam \rdata_comb[30]~227 .sum_lutc_input = "datac";

dffeas \csr_rd_inst_data[31] (
	.clk(clk),
	.d(csr_wrdata[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_rd_inst~combout ),
	.q(\csr_rd_inst_data[31]~q ),
	.prn(vcc));
defparam \csr_rd_inst_data[31] .is_wysiwyg = "true";
defparam \csr_rd_inst_data[31] .power_up = "low";

dffeas \csr_flash_cmd_rd_data_0_data[31] (
	.clk(clk),
	.d(out_rsp_data_31),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_0_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_0_data[31]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_0_data[31] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_0_data[31] .power_up = "low";

dffeas \csr_op_protocol_data[31] (
	.clk(clk),
	.d(csr_wrdata[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_op_protocol~combout ),
	.q(\csr_op_protocol_data[31]~q ),
	.prn(vcc));
defparam \csr_op_protocol_data[31] .is_wysiwyg = "true";
defparam \csr_op_protocol_data[31] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[31]~228 (
	.dataa(avl_csr_address_0),
	.datab(\csr_flash_cmd_rd_data_0_data[31]~q ),
	.datac(avl_csr_address_3),
	.datad(\csr_op_protocol_data[31]~q ),
	.cin(gnd),
	.combout(\rdata_comb[31]~228_combout ),
	.cout());
defparam \rdata_comb[31]~228 .lut_mask = 16'hE5E0;
defparam \rdata_comb[31]~228 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_rd_data_1_data[31] (
	.clk(clk),
	.d(out_rsp_data_31),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\csr_flash_cmd_rd_data_1_data[0]~0_combout ),
	.q(\csr_flash_cmd_rd_data_1_data[31]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_rd_data_1_data[31] .is_wysiwyg = "true";
defparam \csr_flash_cmd_rd_data_1_data[31] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[31]~229 (
	.dataa(\csr_rd_inst_data[31]~q ),
	.datab(avl_csr_address_0),
	.datac(\rdata_comb[31]~228_combout ),
	.datad(\csr_flash_cmd_rd_data_1_data[31]~q ),
	.cin(gnd),
	.combout(\rdata_comb[31]~229_combout ),
	.cout());
defparam \rdata_comb[31]~229 .lut_mask = 16'hF838;
defparam \rdata_comb[31]~229 .sum_lutc_input = "datac";

dffeas \csr_control_data[31] (
	.clk(clk),
	.d(csr_wrdata[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_control~combout ),
	.q(\csr_control_data[31]~q ),
	.prn(vcc));
defparam \csr_control_data[31] .is_wysiwyg = "true";
defparam \csr_control_data[31] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[31]~230 (
	.dataa(\avl_rddata_local[13]~9_combout ),
	.datab(\rdata_comb[31]~229_combout ),
	.datac(\avl_rddata_local[13]~8_combout ),
	.datad(\csr_control_data[31]~q ),
	.cin(gnd),
	.combout(\rdata_comb[31]~230_combout ),
	.cout());
defparam \rdata_comb[31]~230 .lut_mask = 16'hE5E0;
defparam \rdata_comb[31]~230 .sum_lutc_input = "datac";

dffeas \csr_flash_cmd_setting_data[31] (
	.clk(clk),
	.d(csr_wrdata[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_flash_cmd_setting~combout ),
	.q(\csr_flash_cmd_setting_data[31]~q ),
	.prn(vcc));
defparam \csr_flash_cmd_setting_data[31] .is_wysiwyg = "true";
defparam \csr_flash_cmd_setting_data[31] .power_up = "low";

dffeas \csr_wr_inst_data[31] (
	.clk(clk),
	.d(csr_wrdata[31]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_csr_wr_inst~combout ),
	.q(\csr_wr_inst_data[31]~q ),
	.prn(vcc));
defparam \csr_wr_inst_data[31] .is_wysiwyg = "true";
defparam \csr_wr_inst_data[31] .power_up = "low";

cycloneive_lcell_comb \rdata_comb[31]~231 (
	.dataa(avl_csr_address_3),
	.datab(\csr_flash_cmd_setting_data[31]~q ),
	.datac(avl_csr_address_0),
	.datad(\csr_wr_inst_data[31]~q ),
	.cin(gnd),
	.combout(\rdata_comb[31]~231_combout ),
	.cout());
defparam \rdata_comb[31]~231 .lut_mask = 16'hE5E0;
defparam \rdata_comb[31]~231 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[31]~232 (
	.dataa(csr_flash_cmd_wr_data_0_data_31),
	.datab(avl_csr_address_3),
	.datac(\rdata_comb[31]~231_combout ),
	.datad(csr_flash_cmd_wr_data_1_data_31),
	.cin(gnd),
	.combout(\rdata_comb[31]~232_combout ),
	.cout());
defparam \rdata_comb[31]~232 .lut_mask = 16'hF838;
defparam \rdata_comb[31]~232 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[31]~233 (
	.dataa(csr_flash_cmd_addr_data_31),
	.datab(\avl_rddata_local[13]~9_combout ),
	.datac(\rdata_comb[31]~230_combout ),
	.datad(\rdata_comb[31]~232_combout ),
	.cin(gnd),
	.combout(\rdata_comb[31]~233_combout ),
	.cout());
defparam \rdata_comb[31]~233 .lut_mask = 16'hF838;
defparam \rdata_comb[31]~233 .sum_lutc_input = "datac";

cycloneive_lcell_comb \rdata_comb[31]~234 (
	.dataa(\rdata_comb[31]~233_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\avl_rddata_local[13]~10_combout ),
	.cin(gnd),
	.combout(\rdata_comb[31]~234_combout ),
	.cout());
defparam \rdata_comb[31]~234 .lut_mask = 16'h00AA;
defparam \rdata_comb[31]~234 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector32~0 (
	.dataa(stateST_SEND_DUMMY_RSP),
	.datab(out_valid),
	.datac(out_endofpacket),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector32~0_combout ),
	.cout());
defparam \Selector32~0 .lut_mask = 16'hEAEA;
defparam \Selector32~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_csr_flash_cmd_control~0 (
	.dataa(csr_wrdata[0]),
	.datab(csr_wrdata[1]),
	.datac(csr_wrdata[2]),
	.datad(csr_wrdata[3]),
	.cin(gnd),
	.combout(\wr_csr_flash_cmd_control~0_combout ),
	.cout());
defparam \wr_csr_flash_cmd_control~0 .lut_mask = 16'h0002;
defparam \wr_csr_flash_cmd_control~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_csr_flash_cmd_control~1 (
	.dataa(avl_csr_address_1),
	.datab(avl_csr_address_0),
	.datac(csr_wrdata[4]),
	.datad(csr_wrdata[5]),
	.cin(gnd),
	.combout(\wr_csr_flash_cmd_control~1_combout ),
	.cout());
defparam \wr_csr_flash_cmd_control~1 .lut_mask = 16'h0001;
defparam \wr_csr_flash_cmd_control~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_csr_flash_cmd_control~2 (
	.dataa(csr_wrdata[6]),
	.datab(csr_wrdata[7]),
	.datac(csr_wrdata[8]),
	.datad(csr_wrdata[9]),
	.cin(gnd),
	.combout(\wr_csr_flash_cmd_control~2_combout ),
	.cout());
defparam \wr_csr_flash_cmd_control~2 .lut_mask = 16'h0001;
defparam \wr_csr_flash_cmd_control~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_csr_flash_cmd_control~3 (
	.dataa(csr_wrdata[10]),
	.datab(csr_wrdata[11]),
	.datac(csr_wrdata[12]),
	.datad(csr_wrdata[13]),
	.cin(gnd),
	.combout(\wr_csr_flash_cmd_control~3_combout ),
	.cout());
defparam \wr_csr_flash_cmd_control~3 .lut_mask = 16'h0001;
defparam \wr_csr_flash_cmd_control~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_csr_flash_cmd_control~4 (
	.dataa(\wr_csr_flash_cmd_control~0_combout ),
	.datab(\wr_csr_flash_cmd_control~1_combout ),
	.datac(\wr_csr_flash_cmd_control~2_combout ),
	.datad(\wr_csr_flash_cmd_control~3_combout ),
	.cin(gnd),
	.combout(\wr_csr_flash_cmd_control~4_combout ),
	.cout());
defparam \wr_csr_flash_cmd_control~4 .lut_mask = 16'h8000;
defparam \wr_csr_flash_cmd_control~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_csr_flash_cmd_control~5 (
	.dataa(avl_csr_address_3),
	.datab(\wr_csr_control~0_combout ),
	.datac(\wr_csr_flash_cmd_control~4_combout ),
	.datad(avl_csr_address_2),
	.cin(gnd),
	.combout(\wr_csr_flash_cmd_control~5_combout ),
	.cout());
defparam \wr_csr_flash_cmd_control~5 .lut_mask = 16'h0080;
defparam \wr_csr_flash_cmd_control~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_csr_flash_cmd_control~6 (
	.dataa(csr_wrdata[14]),
	.datab(csr_wrdata[15]),
	.datac(csr_wrdata[16]),
	.datad(csr_wrdata[17]),
	.cin(gnd),
	.combout(\wr_csr_flash_cmd_control~6_combout ),
	.cout());
defparam \wr_csr_flash_cmd_control~6 .lut_mask = 16'h0001;
defparam \wr_csr_flash_cmd_control~6 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_csr_flash_cmd_control~7 (
	.dataa(csr_wrdata[18]),
	.datab(csr_wrdata[19]),
	.datac(csr_wrdata[20]),
	.datad(csr_wrdata[21]),
	.cin(gnd),
	.combout(\wr_csr_flash_cmd_control~7_combout ),
	.cout());
defparam \wr_csr_flash_cmd_control~7 .lut_mask = 16'h0001;
defparam \wr_csr_flash_cmd_control~7 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_csr_flash_cmd_control~8 (
	.dataa(csr_wrdata[22]),
	.datab(csr_wrdata[23]),
	.datac(csr_wrdata[24]),
	.datad(csr_wrdata[25]),
	.cin(gnd),
	.combout(\wr_csr_flash_cmd_control~8_combout ),
	.cout());
defparam \wr_csr_flash_cmd_control~8 .lut_mask = 16'h0001;
defparam \wr_csr_flash_cmd_control~8 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_csr_flash_cmd_control~9 (
	.dataa(csr_wrdata[26]),
	.datab(csr_wrdata[27]),
	.datac(csr_wrdata[28]),
	.datad(csr_wrdata[29]),
	.cin(gnd),
	.combout(\wr_csr_flash_cmd_control~9_combout ),
	.cout());
defparam \wr_csr_flash_cmd_control~9 .lut_mask = 16'h0001;
defparam \wr_csr_flash_cmd_control~9 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_csr_flash_cmd_control~10 (
	.dataa(\wr_csr_flash_cmd_control~6_combout ),
	.datab(\wr_csr_flash_cmd_control~7_combout ),
	.datac(\wr_csr_flash_cmd_control~8_combout ),
	.datad(\wr_csr_flash_cmd_control~9_combout ),
	.cin(gnd),
	.combout(\wr_csr_flash_cmd_control~10_combout ),
	.cout());
defparam \wr_csr_flash_cmd_control~10 .lut_mask = 16'h8000;
defparam \wr_csr_flash_cmd_control~10 .sum_lutc_input = "datac";

cycloneive_lcell_comb \wr_csr_flash_cmd_control~11 (
	.dataa(\wr_csr_flash_cmd_control~5_combout ),
	.datab(\wr_csr_flash_cmd_control~10_combout ),
	.datac(csr_wrdata[30]),
	.datad(csr_wrdata[31]),
	.cin(gnd),
	.combout(\wr_csr_flash_cmd_control~11_combout ),
	.cout());
defparam \wr_csr_flash_cmd_control~11 .lut_mask = 16'h0008;
defparam \wr_csr_flash_cmd_control~11 .sum_lutc_input = "datac";

dffeas flash_operation_reg(
	.clk(clk),
	.d(\wr_csr_flash_cmd_control~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\flash_operation_reg~q ),
	.prn(vcc));
defparam flash_operation_reg.is_wysiwyg = "true";
defparam flash_operation_reg.power_up = "low";

cycloneive_lcell_comb \Selector32~1 (
	.dataa(\Selector32~0_combout ),
	.datab(sink_ready),
	.datac(\flash_operation_reg~q ),
	.datad(stateST_IDLE),
	.cin(gnd),
	.combout(\Selector32~1_combout ),
	.cout());
defparam \Selector32~1 .lut_mask = 16'h7770;
defparam \Selector32~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \avl_rddatavalid_local~0 (
	.dataa(hold_waitrequest),
	.datab(avl_csr_read),
	.datac(\flash_operation_reg~q ),
	.datad(stateST_IDLE),
	.cin(gnd),
	.combout(\avl_rddatavalid_local~0_combout ),
	.cout());
defparam \avl_rddatavalid_local~0 .lut_mask = 16'h0008;
defparam \avl_rddatavalid_local~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \csr_rd_inst_data[0]~0 (
	.dataa(csr_wrdata[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\csr_rd_inst_data[0]~0_combout ),
	.cout());
defparam \csr_rd_inst_data[0]~0 .lut_mask = 16'h5555;
defparam \csr_rd_inst_data[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb wr_csr_flash_cmd_wr_data_0(
	.dataa(avl_csr_address_1),
	.datab(avl_csr_address_3),
	.datac(\wr_csr_control~1_combout ),
	.datad(avl_csr_address_0),
	.cin(gnd),
	.combout(\wr_csr_flash_cmd_wr_data_0~combout ),
	.cout());
defparam wr_csr_flash_cmd_wr_data_0.lut_mask = 16'h0080;
defparam wr_csr_flash_cmd_wr_data_0.sum_lutc_input = "datac";

cycloneive_lcell_comb wr_csr_flash_cmd_addr(
	.dataa(avl_csr_address_3),
	.datab(\wr_csr_flash_cmd_addr~0_combout ),
	.datac(\wr_csr_control~0_combout ),
	.datad(avl_csr_address_2),
	.cin(gnd),
	.combout(\wr_csr_flash_cmd_addr~combout ),
	.cout());
defparam wr_csr_flash_cmd_addr.lut_mask = 16'h0080;
defparam wr_csr_flash_cmd_addr.sum_lutc_input = "datac";

cycloneive_lcell_comb wr_csr_flash_cmd_wr_data_1(
	.dataa(avl_csr_address_1),
	.datab(avl_csr_address_0),
	.datac(avl_csr_address_3),
	.datad(\wr_csr_control~1_combout ),
	.cin(gnd),
	.combout(\wr_csr_flash_cmd_wr_data_1~combout ),
	.cout());
defparam wr_csr_flash_cmd_wr_data_1.lut_mask = 16'h8000;
defparam wr_csr_flash_cmd_wr_data_1.sum_lutc_input = "datac";

cycloneive_lcell_comb wr_csr_delay_setting(
	.dataa(avl_csr_address_1),
	.datab(\wr_csr_control~1_combout ),
	.datac(avl_csr_address_0),
	.datad(avl_csr_address_3),
	.cin(gnd),
	.combout(\wr_csr_delay_setting~combout ),
	.cout());
defparam wr_csr_delay_setting.lut_mask = 16'h0008;
defparam wr_csr_delay_setting.sum_lutc_input = "datac";

cycloneive_lcell_comb \csr_clk_baud_rate_data[4]~2 (
	.dataa(csr_wrdata[0]),
	.datab(csr_wrdata[1]),
	.datac(csr_wrdata[2]),
	.datad(csr_wrdata[3]),
	.cin(gnd),
	.combout(\csr_clk_baud_rate_data[4]~2_combout ),
	.cout());
defparam \csr_clk_baud_rate_data[4]~2 .lut_mask = 16'h0001;
defparam \csr_clk_baud_rate_data[4]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \csr_clk_baud_rate_data[4]~4 (
	.dataa(avl_csr_address_0),
	.datab(avl_csr_address_1),
	.datac(csr_wrdata[4]),
	.datad(\csr_clk_baud_rate_data[4]~2_combout ),
	.cin(gnd),
	.combout(\csr_clk_baud_rate_data[4]~4_combout ),
	.cout());
defparam \csr_clk_baud_rate_data[4]~4 .lut_mask = 16'h2002;
defparam \csr_clk_baud_rate_data[4]~4 .sum_lutc_input = "datac";

cycloneive_lcell_comb \csr_clk_baud_rate_data[4]~3 (
	.dataa(\wr_csr_control~0_combout ),
	.datab(\csr_clk_baud_rate_data[4]~4_combout ),
	.datac(avl_csr_address_2),
	.datad(avl_csr_address_3),
	.cin(gnd),
	.combout(\csr_clk_baud_rate_data[4]~3_combout ),
	.cout());
defparam \csr_clk_baud_rate_data[4]~3 .lut_mask = 16'h0008;
defparam \csr_clk_baud_rate_data[4]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \csr_control_data[0]~0 (
	.dataa(csr_wrdata[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\csr_control_data[0]~0_combout ),
	.cout());
defparam \csr_control_data[0]~0 .lut_mask = 16'h5555;
defparam \csr_control_data[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb wr_csr_rd_capturing(
	.dataa(avl_csr_address_1),
	.datab(avl_csr_address_0),
	.datac(\wr_csr_control~1_combout ),
	.datad(avl_csr_address_3),
	.cin(gnd),
	.combout(\wr_csr_rd_capturing~combout ),
	.cout());
defparam wr_csr_rd_capturing.lut_mask = 16'h0080;
defparam wr_csr_rd_capturing.sum_lutc_input = "datac";

cycloneive_lcell_comb \csr_wr_inst_data[1]~0 (
	.dataa(csr_wrdata[1]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\csr_wr_inst_data[1]~0_combout ),
	.cout());
defparam \csr_wr_inst_data[1]~0 .lut_mask = 16'h5555;
defparam \csr_wr_inst_data[1]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \csr_rd_inst_data[1]~1 (
	.dataa(csr_wrdata[1]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\csr_rd_inst_data[1]~1_combout ),
	.cout());
defparam \csr_rd_inst_data[1]~1 .lut_mask = 16'h5555;
defparam \csr_rd_inst_data[1]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \csr_clk_baud_rate_data[4]~5 (
	.dataa(csr_wrdata[4]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\csr_clk_baud_rate_data[4]~5_combout ),
	.cout());
defparam \csr_clk_baud_rate_data[4]~5 .lut_mask = 16'h5555;
defparam \csr_clk_baud_rate_data[4]~5 .sum_lutc_input = "datac";

cycloneive_lcell_comb \csr_wr_inst_data[12]~1 (
	.dataa(csr_wrdata[12]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\csr_wr_inst_data[12]~1_combout ),
	.cout());
defparam \csr_wr_inst_data[12]~1 .lut_mask = 16'h5555;
defparam \csr_wr_inst_data[12]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \csr_wr_inst_data[13]~2 (
	.dataa(csr_wrdata[13]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\csr_wr_inst_data[13]~2_combout ),
	.cout());
defparam \csr_wr_inst_data[13]~2 .lut_mask = 16'h5555;
defparam \csr_wr_inst_data[13]~2 .sum_lutc_input = "datac";

cycloneive_lcell_comb \csr_wr_inst_data[14]~3 (
	.dataa(csr_wrdata[14]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\csr_wr_inst_data[14]~3_combout ),
	.cout());
defparam \csr_wr_inst_data[14]~3 .lut_mask = 16'h5555;
defparam \csr_wr_inst_data[14]~3 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector36~0 (
	.dataa(saved_grant_1),
	.datab(stateST_SEND_DATA_1),
	.datac(src_payload_0),
	.datad(Selector18),
	.cin(gnd),
	.combout(\Selector36~0_combout ),
	.cout());
defparam \Selector36~0 .lut_mask = 16'hA800;
defparam \Selector36~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector36~1 (
	.dataa(\Selector32~0_combout ),
	.datab(in_cmd_channel_reg_1),
	.datac(stateST_WAIT_RSP),
	.datad(\Selector36~0_combout ),
	.cin(gnd),
	.combout(\Selector36~1_combout ),
	.cout());
defparam \Selector36~1 .lut_mask = 16'hFF70;
defparam \Selector36~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector33~0 (
	.dataa(\flash_operation_reg~q ),
	.datab(stateST_SEND_HEADER),
	.datac(stateST_IDLE),
	.datad(sink1_ready),
	.cin(gnd),
	.combout(\Selector33~0_combout ),
	.cout());
defparam \Selector33~0 .lut_mask = 16'h0ACE;
defparam \Selector33~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Selector35~0 (
	.dataa(more_than_4bytes_data1),
	.datab(stateST_SEND_DATA_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector35~0_combout ),
	.cout());
defparam \Selector35~0 .lut_mask = 16'h8888;
defparam \Selector35~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal16~0 (
	.dataa(\csr_flash_cmd_setting_data[12]~q ),
	.datab(\csr_flash_cmd_setting_data[13]~q ),
	.datac(\csr_flash_cmd_setting_data[14]~q ),
	.datad(\csr_flash_cmd_setting_data[15]~q ),
	.cin(gnd),
	.combout(\Equal16~0_combout ),
	.cout());
defparam \Equal16~0 .lut_mask = 16'h0002;
defparam \Equal16~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \has_data_in~0 (
	.dataa(\Equal16~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\csr_flash_cmd_setting_data[11]~q ),
	.cin(gnd),
	.combout(\has_data_in~0_combout ),
	.cout());
defparam \has_data_in~0 .lut_mask = 16'h5500;
defparam \has_data_in~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \LessThan0~0 (
	.dataa(\csr_flash_cmd_setting_data[15]~q ),
	.datab(\csr_flash_cmd_setting_data[14]~q ),
	.datac(\csr_flash_cmd_setting_data[13]~q ),
	.datad(\csr_flash_cmd_setting_data[12]~q ),
	.cin(gnd),
	.combout(\LessThan0~0_combout ),
	.cout());
defparam \LessThan0~0 .lut_mask = 16'hEAEE;
defparam \LessThan0~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \has_data_out~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\csr_flash_cmd_setting_data[11]~q ),
	.datad(\Equal16~0_combout ),
	.cin(gnd),
	.combout(\has_data_out~0_combout ),
	.cout());
defparam \has_data_out~0 .lut_mask = 16'h000F;
defparam \has_data_out~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \numb_data[0]~0 (
	.dataa(\csr_flash_cmd_setting_data[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\numb_data[0]~0_combout ),
	.cout());
defparam \numb_data[0]~0 .lut_mask = 16'h5555;
defparam \numb_data[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal13~0 (
	.dataa(gnd),
	.datab(\csr_flash_cmd_setting_data[8]~q ),
	.datac(\csr_flash_cmd_setting_data[9]~q ),
	.datad(\csr_flash_cmd_setting_data[10]~q ),
	.cin(gnd),
	.combout(\Equal13~0_combout ),
	.cout());
defparam \Equal13~0 .lut_mask = 16'hFFFC;
defparam \Equal13~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal14~0 (
	.dataa(\csr_flash_cmd_setting_data[10]~q ),
	.datab(gnd),
	.datac(\csr_flash_cmd_setting_data[8]~q ),
	.datad(\csr_flash_cmd_setting_data[9]~q ),
	.cin(gnd),
	.combout(\Equal14~0_combout ),
	.cout());
defparam \Equal14~0 .lut_mask = 16'h000A;
defparam \Equal14~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \opcode[0]~0 (
	.dataa(\csr_flash_cmd_setting_data[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\opcode[0]~0_combout ),
	.cout());
defparam \opcode[0]~0 .lut_mask = 16'h5555;
defparam \opcode[0]~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \opcode[2]~1 (
	.dataa(\csr_flash_cmd_setting_data[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\opcode[2]~1_combout ),
	.cout());
defparam \opcode[2]~1 .lut_mask = 16'h5555;
defparam \opcode[2]~1 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal15~0 (
	.dataa(\csr_flash_cmd_setting_data[17]~q ),
	.datab(\csr_flash_cmd_setting_data[18]~q ),
	.datac(\csr_flash_cmd_setting_data[19]~q ),
	.datad(\csr_flash_cmd_setting_data[20]~q ),
	.cin(gnd),
	.combout(\Equal15~0_combout ),
	.cout());
defparam \Equal15~0 .lut_mask = 16'h0001;
defparam \Equal15~0 .sum_lutc_input = "datac";

cycloneive_lcell_comb \Equal15~1 (
	.dataa(\Equal15~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\csr_flash_cmd_setting_data[16]~q ),
	.cin(gnd),
	.combout(\Equal15~1_combout ),
	.cout());
defparam \Equal15~1 .lut_mask = 16'hFF55;
defparam \Equal15~1 .sum_lutc_input = "datac";

endmodule

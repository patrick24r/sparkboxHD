module engineTop(
	input clk, 
	input reset, 
	input cmd, 
	input cmdData, 
	input flashData, 
	input ramData, 
	output fontIndex, 
	output fontSize, 
	output ramAddr, 
	output [4:0] layer, 
	output [5:0] paletteIndex, 
	output frameDone);
	
	
endmodule
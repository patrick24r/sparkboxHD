// qspi_inf_mux.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module qspi_inf_mux (
		input  wire        clk,                 //       clk.clk
		input  wire        reset,               // clk_reset.reset
		input  wire        src_ready,           //       src.ready
		output wire        src_valid,           //          .valid
		output wire [3:0]  src_data,            //          .data
		output wire [11:0] src_channel,         //          .channel
		output wire        src_startofpacket,   //          .startofpacket
		output wire        src_endofpacket,     //          .endofpacket
		output wire        sink0_ready,         //     sink0.ready
		input  wire        sink0_valid,         //          .valid
		input  wire [11:0] sink0_channel,       //          .channel
		input  wire [3:0]  sink0_data,          //          .data
		input  wire        sink0_startofpacket, //          .startofpacket
		input  wire        sink0_endofpacket,   //          .endofpacket
		output wire        sink1_ready,         //     sink1.ready
		input  wire        sink1_valid,         //          .valid
		input  wire [11:0] sink1_channel,       //          .channel
		input  wire [3:0]  sink1_data,          //          .data
		input  wire        sink1_startofpacket, //          .startofpacket
		input  wire        sink1_endofpacket,   //          .endofpacket
		output wire        sink2_ready,         //     sink2.ready
		input  wire        sink2_valid,         //          .valid
		input  wire [11:0] sink2_channel,       //          .channel
		input  wire [3:0]  sink2_data,          //          .data
		input  wire        sink2_startofpacket, //          .startofpacket
		input  wire        sink2_endofpacket    //          .endofpacket
	);

	flashLoader_intel_generic_serial_flash_interface_top_0_qspi_inf_inst_qspi_inf_mux_qspi_inf_mux qspi_inf_mux (
		.clk                 (clk),                 //       clk.clk
		.reset               (reset),               // clk_reset.reset
		.src_ready           (src_ready),           //       src.ready
		.src_valid           (src_valid),           //          .valid
		.src_data            (src_data),            //          .data
		.src_channel         (src_channel),         //          .channel
		.src_startofpacket   (src_startofpacket),   //          .startofpacket
		.src_endofpacket     (src_endofpacket),     //          .endofpacket
		.sink0_ready         (sink0_ready),         //     sink0.ready
		.sink0_valid         (sink0_valid),         //          .valid
		.sink0_channel       (sink0_channel),       //          .channel
		.sink0_data          (sink0_data),          //          .data
		.sink0_startofpacket (sink0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (sink0_endofpacket),   //          .endofpacket
		.sink1_ready         (sink1_ready),         //     sink1.ready
		.sink1_valid         (sink1_valid),         //          .valid
		.sink1_channel       (sink1_channel),       //          .channel
		.sink1_data          (sink1_data),          //          .data
		.sink1_startofpacket (sink1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (sink1_endofpacket),   //          .endofpacket
		.sink2_ready         (sink2_ready),         //     sink2.ready
		.sink2_valid         (sink2_valid),         //          .valid
		.sink2_channel       (sink2_channel),       //          .channel
		.sink2_data          (sink2_data),          //          .data
		.sink2_startofpacket (sink2_startofpacket), //          .startofpacket
		.sink2_endofpacket   (sink2_endofpacket)    //          .endofpacket
	);

endmodule

module controllerTop(

);

endmodule
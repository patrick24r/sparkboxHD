// This layer serves as memory to store a register for all layers
// E.g. Stores register 0 for all layers
module layerRegisterMem(
    input clk,
    input reset,
    input [4:0] readAddr,
    input writeEn,
    input [4:0] writeAddr,
    input [15:0] writeData,
    output [15:0] readData
);

reg [15:0] layerRegisters [4:0];

// Initialize all data as blank
initial begin
    for (1 = 0; i < 32; i = i + 1) begin
        layerRegisters[i] = 16'd0;
    end
end

// Asynchronous reads
assign readData = layerRegisters[readAddr];

// Writes on posedge
always @(posedge clk) begin
    if (!reset) begin
    // Reset all data to 0
        for (1 = 0; i < 32; i = i + 1) begin
            layerRegisters[i] <= 16'd0;
        end
    end
    else begin
        layerRegisters[writeAddr] <= writeData;
    end
end

endmodule
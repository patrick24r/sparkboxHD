// flashLoader.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module flashLoader (
		input  wire [5:0]  avl_csr_address,       // avl_csr.address
		input  wire        avl_csr_read,          //        .read
		output wire [31:0] avl_csr_readdata,      //        .readdata
		input  wire        avl_csr_write,         //        .write
		input  wire [31:0] avl_csr_writedata,     //        .writedata
		output wire        avl_csr_waitrequest,   //        .waitrequest
		output wire        avl_csr_readdatavalid, //        .readdatavalid
		input  wire        avl_mem_write,         // avl_mem.write
		input  wire [6:0]  avl_mem_burstcount,    //        .burstcount
		output wire        avl_mem_waitrequest,   //        .waitrequest
		input  wire        avl_mem_read,          //        .read
		input  wire [20:0] avl_mem_address,       //        .address
		input  wire [31:0] avl_mem_writedata,     //        .writedata
		output wire [31:0] avl_mem_readdata,      //        .readdata
		output wire        avl_mem_readdatavalid, //        .readdatavalid
		input  wire [3:0]  avl_mem_byteenable,    //        .byteenable
		input  wire        clk_clk,               //     clk.clk
		input  wire        reset_reset            //   reset.reset
	);

	flashLoader_intel_generic_serial_flash_interface_top_0 #(
		.DEVICE_FAMILY ("Cyclone IV E"),
		.CHIP_SELS     (1)
	) intel_generic_serial_flash_interface_top_0 (
		.avl_csr_address       (avl_csr_address),       // avl_csr.address
		.avl_csr_read          (avl_csr_read),          //        .read
		.avl_csr_readdata      (avl_csr_readdata),      //        .readdata
		.avl_csr_write         (avl_csr_write),         //        .write
		.avl_csr_writedata     (avl_csr_writedata),     //        .writedata
		.avl_csr_waitrequest   (avl_csr_waitrequest),   //        .waitrequest
		.avl_csr_readdatavalid (avl_csr_readdatavalid), //        .readdatavalid
		.avl_mem_write         (avl_mem_write),         // avl_mem.write
		.avl_mem_burstcount    (avl_mem_burstcount),    //        .burstcount
		.avl_mem_waitrequest   (avl_mem_waitrequest),   //        .waitrequest
		.avl_mem_read          (avl_mem_read),          //        .read
		.avl_mem_address       (avl_mem_address),       //        .address
		.avl_mem_writedata     (avl_mem_writedata),     //        .writedata
		.avl_mem_readdata      (avl_mem_readdata),      //        .readdata
		.avl_mem_readdatavalid (avl_mem_readdatavalid), //        .readdatavalid
		.avl_mem_byteenable    (avl_mem_byteenable),    //        .byteenable
		.clk_clk               (clk_clk),               //     clk.clk
		.reset_reset           (reset_reset)            //   reset.reset
	);

endmodule

module simLcdTester(
);
endmodule